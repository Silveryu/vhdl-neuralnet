----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 05/31/2018 02:49:06 PM
-- Design Name: 
-- Module Name: weight_unit_tb - Stimulus
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;


library work;
use work.custom_type.all;


entity mat_mult_tb is
end mat_mult_tb;

architecture Stimulus of mat_mult_tb is

    constant TIME_DELTA: time := 10 ns; -- clock wait time in ns
    constant N : positive := 784;
    constant M : positive := 2;

    
    signal X : WORD_ARRAY(0 to N-1) := ( X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0030", X"0121", X"0121", X"0121", X"07E8", X"0888", X"0AFA", X"01A2", X"0A6A", X"1000", X"0F80", X"07F8", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"01E2", X"0243", X"05E6", X"09AA", X"0AAA", X"0FE0", X"0FE0", X"0FE0", X"0FE0", X"0FE0", X"0E1E", X"0ACA", X"0FE0", X"0F30", X"0C3C", X"0404", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0313", X"0EEE", X"0FE0", X"0FE0", X"0FE0", X"0FE0", X"0FE0", X"0FE0", X"0FE0", X"0FE0", X"0FC0", X"05D6", X"0525", X"0525", X"0384", X"0273", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0121", X"0DBE", X"0FE0", X"0FE0", X"0FE0", X"0FE0", X"0FE0", X"0C6C", X"0B6C", X"0F80", X"0F20", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0505", X"09CA", X"06B7", X"0FE0", X"0FE0", X"0CDC", X"00B1", X"0000", X"02B3", X"09AA", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"00E1", X"0010", X"09AA", X"0FE0", X"05A6", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"08B8", X"0FE0", X"0BEC", X"0020", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"00B1", X"0BEC", X"0FE0", X"0464", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0232", X"0F20", X"0E1E", X"0A0A", X"06C7", X"0010", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0515", X"0F10", X"0FE0", X"0FE0", X"0777", X"0192", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"02D3", X"0BAC", X"0FE0", X"0FE0", X"096A", X"01B2", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0101", X"05D6", X"0FD0", X"0FE0", X"0BBC", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0FA0", X"0FE0", X"0FA0", X"0404", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"02E3", X"0828", X"0B7C", X"0FE0", X"0FE0", X"0CFC", X"0020", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0273", X"094A", X"0E5E", X"0FE0", X"0FE0", X"0FE0", X"0FB0", X"0B6C", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0182", X"0727", X"0DDE", X"0FE0", X"0FE0", X"0FE0", X"0FE0", X"0C9C", X"04E5", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0172", X"0424", X"0D5E", X"0FE0", X"0FE0", X"0FE0", X"0FE0", X"0C6C", X"0515", X"0020", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0121", X"0ABA", X"0DBE", X"0FE0", X"0FE0", X"0FE0", X"0FE0", X"0C3C", X"0505", X"0091", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0374", X"0ACA", X"0E2E", X"0FE0", X"0FE0", X"0FE0", X"0FE0", X"0F50", X"0858", X"00B1", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0888", X"0FE0", X"0FE0", X"0FE0", X"0D4E", X"0878", X"0848", X"0101", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000");
    signal Z : WORD_ARRAY(0 to M-1);
    
    signal W1 : WORD_MAT(0 to M-1, 0 to N-1) := (	
        (X"FFA8", X"FF30", X"FEFF", X"FEBA", X"FFF9", X"FFE1", X"FF24", X"0021", X"005F", X"FF24", X"0081", X"FFEC", X"FFBD", X"00B6", X"FF8F", X"FFFB", X"0082", X"FF31", X"00B3", X"FECA", X"022D", X"003A", X"0060", X"FFA9", X"0007", X"0069", X"FF74", X"02A6", X"FEEB", X"003C", X"015D", X"00CC", X"0063", X"0045", X"FF00", X"006D", X"0069", X"FF2D", X"FE47", X"FFF8", X"FFD2", X"0170", X"FE4E", X"0061", X"009F", X"01AA", X"FDD1", X"FE3D", X"FE38", X"004B", X"FF75", X"FF90", X"001C", X"FF07", X"FE7F", X"01AF", X"FF15", X"FE91", X"0035", X"0125", X"FF1D", X"FF4F", X"FEFE", X"FFE8", X"FEEC", X"FE3E", X"FAAB", X"FC43", X"FB25", X"FDE2", X"F9A2", X"FB22", X"FCC9", X"FC84", X"FC0F", X"FE45", X"FAC1", X"FACC", X"FAA9", X"FD40", X"FE28", X"01D2", X"FF4A", X"00EE", X"FF22", X"FE77", X"FEDD", X"0042", X"FEFE", X"FE0B", X"FD8D", X"FD2F", X"FDB2", X"FCB1", X"F9AC", X"FA53", X"FA04", X"FB05", X"FB4B", X"FBDD", X"FB60", X"FC9E", X"F950", X"F952", X"FA0E", X"FB86", X"FD6A", X"FDC4", X"FE63", X"FE50", X"FEE7", X"FFE7", X"015F", X"0027", X"0007", X"00B3", X"FD52", X"FBDF", X"FBED", X"FBB3", X"F74F", X"F93E", X"F83D", X"FAA1", X"F9A8", X"F9BB", X"FAD5", X"FC30", X"F750", X"F8AB", X"F92D", X"F807", X"F97D", X"FB67", X"FDBE", X"FE44", X"FF5B", X"FEAF", X"01A3", X"FE7C", X"009B", X"FFB4", X"FF2D", X"FF31", X"FD78", X"FB8E", X"FBBC", X"FA09", X"F96F", X"FB21", X"FBDB", X"FD9A", X"FDD9", X"FD92", X"FBB8", X"F812", X"F6B7", X"F7DF", X"F939", X"FBF0", X"FD68", X"FF59", X"FF6B", X"FB83", X"FDE9", X"003E", X"FFFB", X"FE47", X"FF0B", X"FE7C", X"0157", X"FFC1", X"00E2", X"FF58", X"FD23", X"FB4A", X"FB8A", X"F92C", X"FD15", X"FDEF", X"FDC6", X"FFB0", X"0185", X"023E", X"03EC", X"02A0", X"0287", X"0218", X"0076", X"0183", X"0038", X"FF65", X"FF89", X"01F1", X"00A7", X"FE3B", X"FFB3", X"FEBF", X"00E8", X"FF09", X"FC8F", X"FA33", X"FAF3", X"FBD4", X"FBD7", X"FC6C", X"FFD0", X"0172", X"0330", X"055C", X"04F9", X"082D", X"0891", X"06F9", X"0646", X"03E4", X"0270", X"0245", X"FF0E", X"00E3", X"0600", X"087F", X"01A1", X"FDBB", X"0245", X"022D", X"FEC6", X"FCBB", X"F86F", X"FABE", X"FB2E", X"FE27", X"FF87", X"FF24", X"0073", X"0282", X"030C", X"0585", X"0562", X"05E6", X"0820", X"0527", X"05B1", X"0318", X"0143", X"FFBE", X"FF99", X"07F7", X"0C52", X"0C17", X"0488", X"00A6", X"0051", X"03BD", X"FF9C", X"FE79", X"FA4A", X"FE40", X"FF85", X"FF0D", X"FE67", X"0011", X"00F9", X"0190", X"01AB", X"0540", X"0680", X"04D1", X"039C", X"049A", X"0526", X"01BC", X"00BD", X"FF83", X"028C", X"08E7", X"0D6A", X"0C88", X"0665", X"02E8", X"0188", X"030E", X"02A3", X"FE35", X"FF1F", X"0134", X"01E9", X"00A3", X"0128", X"01B6", X"029E", X"03C6", X"0367", X"04F8", X"0554", X"0191", X"0310", X"00B4", X"0234", X"FFA0", X"0152", X"0301", X"050D", X"0917", X"0BB8", X"0A62", X"06BB", X"02D0", X"0027", X"02DE", X"019B", X"007D", X"016E", X"0393", X"0461", X"02C2", X"034C", X"01F9", X"004D", X"0390", X"036F", X"0342", X"01A4", X"FF12", X"FDE8", X"0091", X"0186", X"00B2", X"02F7", X"0551", X"053A", X"04F4", X"062E", X"0746", X"0509", X"0020", X"0074", X"02D7", X"0481", X"059A", X"0549", X"07C3", X"0617", X"0287", X"005D", X"005C", X"020E", X"0137", X"01B8", X"FFCC", X"FE8D", X"FC7E", X"FA8D", X"FD74", X"0037", X"02BF", X"04DB", X"03B9", X"04F8", X"02A4", X"FDE4", X"FF48", X"00BD", X"034F", X"FFE7", X"029B", X"039E", X"03A6", X"084C", X"066E", X"03B1", X"04DA", X"0152", X"00F7", X"013B", X"0002", X"FFD9", X"FC34", X"FD8D", X"FCED", X"FAA8", X"FCDA", X"FCC2", X"001D", X"0365", X"0088", X"009C", X"FEF7", X"FF59", X"FEA9", X"FD19", X"FF0F", X"0173", X"0047", X"03F8", X"0026", X"0136", X"01A0", X"0269", X"0144", X"0026", X"0060", X"0323", X"FFAF", X"FCF5", X"FC08", X"FAE0", X"F9EB", X"FBD1", X"FD4F", X"FD8F", X"FE0E", X"FFCC", X"FFCA", X"FFFE", X"0082", X"01A2", X"FD1A", X"0084", X"00A0", X"025F", X"FFC5", X"F991", X"FB9A", X"FF89", X"0150", X"FEFC", X"FFD6", X"FE3D", X"0077", X"02E9", X"FE98", X"FC47", X"F9EA", X"F905", X"FC5A", X"FB77", X"FF6A", X"FE58", X"FCE9", X"FEB7", X"FDB7", X"FE61", X"FE9B", X"0298", X"FD4C", X"FC2E", X"FF13", X"FF48", X"FE82", X"FAEB", X"FA20", X"FE72", X"FF2C", X"0031", X"FE7C", X"FEAE", X"FDDD", X"012E", X"0006", X"FB87", X"F840", X"F864", X"FB4D", X"FC71", X"00EE", X"FB84", X"FC7C", X"FBBC", X"FCF3", X"FCC7", X"FC14", X"FF11", X"FC8D", X"FA18", X"FD3D", X"FEC4", X"FEC7", X"F8EB", X"FB45", X"FE30", X"01FD", X"0180", X"FE5E", X"FFD4", X"012E", X"02D6", X"FF92", X"FB77", X"FAA7", X"FC2E", X"FDB5", X"FE4D", X"FE6B", X"FCCA", X"FA49", X"FD38", X"FCF9", X"FCAD", X"FB50", X"FEE1", X"FD58", X"FBAF", X"024C", X"041B", X"FF21", X"FAE3", X"F75D", X"FE7E", X"0133", X"00B8", X"005D", X"0156", X"01E9", X"0216", X"01EC", X"FDB4", X"FE19", X"FED6", X"0045", X"FCF8", X"FDF9", X"FC22", X"FD9F", X"FF20", X"FCF9", X"FF81", X"FD3E", X"FB94", X"FBB7", X"FB8C", X"FB19", X"009E", X"02D8", X"00D0", X"F63F", X"FE6D", X"FE7C", X"0074", X"01CA", X"03D3", X"0151", X"0166", X"0022", X"00F1", X"0032", X"FDD0", X"FCDE", X"FC09", X"FC16", X"FD57", X"FCF7", X"FEF0", X"FCA4", X"FD29", X"FDE3", X"007F", X"FD35", X"FBA6", X"FFD6", X"002F", X"0027", X"FDD7", X"FA4F", X"FDBD", X"0008", X"00D8", X"008D", X"00CE", X"00C0", X"001C", X"FE72", X"FF2F", X"005B", X"FC53", X"FB78", X"FB69", X"FBF7", X"FB52", X"FC8B", X"FC71", X"FBDE", X"FD66", X"FC8E", X"005B", X"0122", X"FCCD", X"012E", X"000A", X"FE2B", X"FA83", X"FBAC", X"FFBD", X"01F7", X"0078", X"018A", X"0127", X"00A5", X"00A0", X"FE98", X"FD65", X"FC0C", X"FAF8", X"FA72", X"FB52", X"FC74", X"F9CC", X"FA8B", X"FD97", X"FB16", X"FCC3", X"FC24", X"018E", X"01A8", X"FE7E", X"003E", X"00F3", X"FEAE", X"F998", X"F993", X"FDCA", X"FD50", X"00F7", X"01CC", X"0323", X"008D", X"0110", X"FF93", X"01C6", X"FECA", X"FF3C", X"FCC4", X"FD44", X"FD15", X"FC72", X"FC18", X"FBF1", X"FAE0", X"FE37", X"00A8", X"0269", X"0181", X"FD7E", X"00DB", X"FFC9", X"015F", X"FAFB", X"F98E", X"F9FF", X"FE14", X"0009", X"0074", X"0154", X"01B1", X"018C", X"02D1", X"0001", X"FFC6", X"FFE9", X"0058", X"FEF8", X"FD63", X"FB62", X"FAAC", X"FDD4", X"FBF0", X"00E4", X"0571", X"0435", X"FF8C", X"FB99", X"002F", X"00BD", X"FF74", X"FEC2", X"0037", X"FFB0", X"02B2", X"022E", X"0060", X"FF87", X"FE22", X"FE61", X"0061", X"01DB", X"029B", X"00A0", X"0196", X"00F4", X"0343", X"0275", X"00A9", X"02E5", X"016B", X"0266", X"04A9", X"01A3", X"FD83", X"FD97", X"000F", X"00E3", X"FFAB", X"FEF9", X"04D1", X"02A2", X"0346", X"008E", X"025F", X"00D3", X"00AE", X"FF3F", X"009A", X"02CD", X"0440", X"0419", X"0678", X"06E3", X"0753", X"07F2", X"0786", X"0740", X"073E", X"041D", X"068C", X"03FF", X"0014", X"FDBB", X"0042", X"FFEA", X"0065", X"FFFD", X"013E", X"029D", X"0405", X"0662", X"04CF", X"05C8", X"0992", X"0A6F", X"0A6E", X"09C7", X"0A30", X"0E98", X"0B3E", X"0963", X"097E", X"07E8", X"087C", X"07FF", X"0877", X"06B3", X"0308", X"00DA", X"FEA0", X"FFC1", X"001E", X"0090", X"FFFB", X"FFA7", X"FFD0", X"018C", X"FF5B", X"0151", X"02D7", X"0448", X"059E", X"0524", X"042B", X"0683", X"0464", X"067E", X"04DD", X"0763", X"0696", X"06CB", X"0331", X"046B", X"03FD", X"03BF", X"0077", X"FF4B", X"003B", X"00ED", X"00E7"),
        (X"FFFD", X"FF64", X"FFD7", X"FFFC", X"0012", X"0026", X"004F", X"0077", X"01A5", X"0019", X"FFA3", X"FFCC", X"FF7E", X"FFA2", X"00BA", X"FFD4", X"FF30", X"FFA7", X"0046", X"00EF", X"00AC", X"FFA9", X"00CE", X"FF38", X"FF39", X"01C1", X"FF80", X"FF43", X"0122", X"00D2", X"FF73", X"FED9", X"0177", X"FF3D", X"FFDA", X"0058", X"0274", X"0268", X"0025", X"FF8F", X"0130", X"00A7", X"FFFB", X"FDF8", X"FBC9", X"FDAD", X"00F5", X"016A", X"0276", X"01A0", X"00CC", X"0014", X"FF6C", X"FFD6", X"FF71", X"00EC", X"FECA", X"0079", X"FF44", X"0009", X"008B", X"015B", X"00A6", X"0283", X"041C", X"01B0", X"01F6", X"008E", X"01D3", X"FF51", X"00E5", X"FD70", X"FD3F", X"FE2D", X"FEB9", X"00E3", X"01D2", X"034F", X"035B", X"02A5", X"030F", X"008F", X"FFF7", X"0096", X"0163", X"FF19", X"FF2C", X"FEFA", X"0002", X"0311", X"04A0", X"0207", X"FFE1", X"FFC0", X"017C", X"021B", X"0187", X"FE7C", X"0144", X"0075", X"000F", X"FFCF", X"0274", X"03E0", X"00E4", X"0264", X"0480", X"039D", X"02D2", X"006F", X"0119", X"0082", X"0022", X"00F1", X"FD88", X"FDF0", X"03A7", X"0403", X"0390", X"0120", X"FE8D", X"FF99", X"FDAE", X"FCB8", X"FD4A", X"FCE7", X"FAB7", X"F8C4", X"FA6A", X"FD1A", X"FB77", X"FD8B", X"FE33", X"FD83", X"0134", X"00F2", X"FE8C", X"FB4D", X"FD67", X"FEA9", X"FFDB", X"FE72", X"FF27", X"FCB3", X"037C", X"027A", X"0344", X"0220", X"045B", X"0128", X"FF17", X"FD3B", X"FC91", X"F9D0", X"FAF2", X"FAED", X"F9CD", X"FA19", X"FBA6", X"FB38", X"F927", X"F769", X"FB63", X"FE4E", X"FCF0", X"FDB8", X"FC99", X"0192", X"012C", X"FF6F", X"FE2B", X"01E5", X"02FD", X"038B", X"0224", X"053F", X"044C", X"0394", X"FEE4", X"FD38", X"FE34", X"FB5C", X"FE27", X"FF2A", X"FEC7", X"FEC2", X"FD27", X"FA6D", X"FBBA", X"FCB2", X"FBA9", X"FB49", X"FC9D", X"FBCA", X"FFF4", X"FD1F", X"0137", X"003B", X"02A8", X"044D", X"01DC", X"02CD", X"0344", X"034F", X"02AB", X"00BC", X"FF42", X"FE97", X"FF30", X"FE79", X"FE0B", X"00D6", X"FED1", X"FED2", X"FB7B", X"FACA", X"FD6E", X"FAAD", X"FBD2", X"FB5A", X"FAF3", X"FD8C", X"FD72", X"FE0B", X"FF6A", X"02DD", X"01C7", X"0180", X"01AF", X"02D7", X"0253", X"0361", X"01E6", X"025D", X"0024", X"FDA3", X"FE2E", X"FE81", X"00E2", X"FE93", X"FCD6", X"FBFE", X"FC69", X"FC02", X"FC8D", X"FB54", X"FB4E", X"F8AF", X"FB83", X"FC81", X"FC4B", X"FBED", X"FF20", X"0427", X"FFC4", X"0191", X"00DC", X"0187", X"01E2", X"01A6", X"0171", X"01F5", X"00E5", X"001B", X"0015", X"0165", X"00E3", X"FE66", X"FC36", X"FA44", X"FD04", X"FD69", X"FCAD", X"FD1C", X"FC16", X"F9F0", X"F8C8", X"F4E0", X"FAED", X"01F6", X"FF36", X"027B", X"FF75", X"00DF", X"0007", X"0144", X"0134", X"01BE", X"034C", X"00C4", X"000F", X"0015", X"01E7", X"0154", X"FEF6", X"FD4A", X"FD02", X"FFF4", X"FFFF", X"FFA8", X"FD07", X"FCF8", X"FBEA", X"F87E", X"F4D3", X"F443", X"F9BD", X"0026", X"0061", X"00D9", X"0354", X"02B0", X"0181", X"0153", X"0106", X"024F", X"035E", X"03D1", X"02F6", X"0289", X"0225", X"FF52", X"FDC5", X"FF15", X"02A1", X"01C4", X"0215", X"FFE5", X"0132", X"00C2", X"FEA1", X"F9DF", X"F387", X"F3C5", X"F7F0", X"FD69", X"01EC", X"01FF", X"04B9", X"0081", X"0354", X"0050", X"016B", X"039E", X"0420", X"0164", X"0240", X"0389", X"FFD6", X"FCB9", X"FC03", X"01D5", X"05B2", X"04AC", X"05F3", X"02DA", X"0247", X"0361", X"04CD", X"0334", X"FA98", X"F82D", X"F93A", X"FE31", X"FF8A", X"FF8F", X"0460", X"FEF7", X"0390", X"030A", X"04F0", X"0321", X"0259", X"0009", X"015B", X"02B0", X"FEE2", X"FCD0", X"FE8D", X"0378", X"05C2", X"046A", X"0402", X"03C1", X"04DB", X"074E", X"081A", X"05D5", X"00C8", X"FD95", X"F89C", X"FCFC", X"FDB5", X"02BA", X"0338", X"017D", X"01BE", X"0188", X"033D", X"02C3", X"0169", X"0019", X"0011", X"00C4", X"FE36", X"FCBF", X"FD86", X"0591", X"0529", X"02B7", X"0448", X"0562", X"0746", X"069F", X"078C", X"04F8", X"02E8", X"01D5", X"F978", X"FE40", X"FFF6", X"00F6", X"022B", X"FF9E", X"0015", X"0023", X"0101", X"02DD", X"0083", X"FCFB", X"FF86", X"01B3", X"0026", X"FD5A", X"0093", X"0582", X"035C", X"050A", X"02DA", X"062A", X"08C7", X"073A", X"0834", X"0454", X"004F", X"FFFC", X"FCA0", X"FDD6", X"0157", X"FF63", X"FF24", X"FC46", X"FC5D", X"FE0F", X"0242", X"02B1", X"013A", X"FD22", X"FF8C", X"002E", X"FF12", X"FF5C", X"035D", X"060F", X"038F", X"0369", X"04B6", X"0487", X"0799", X"0429", X"026F", X"009B", X"FD43", X"FE74", X"FCCA", X"FD68", X"00A0", X"FFEB", X"0031", X"FB93", X"FCFF", X"FBF7", X"FF17", X"01E4", X"0170", X"0027", X"001E", X"03A6", X"018C", X"04DE", X"0483", X"0431", X"0349", X"04E8", X"04A6", X"0266", X"03A4", X"03CB", X"001F", X"FD89", X"FCB5", X"0025", X"FDF1", X"FE76", X"0288", X"0012", X"00EE", X"FE10", X"FCB5", X"FE07", X"FC99", X"FD41", X"FCD9", X"FD1B", X"FF12", X"0208", X"028A", X"0129", X"0153", X"02A2", X"0209", X"00E3", X"FFC8", X"FF55", X"FF42", X"FDF0", X"FC87", X"FC1F", X"F8A8", X"FF98", X"0123", X"FDA3", X"0016", X"FD4E", X"FFD7", X"FC4F", X"FD30", X"FE95", X"FED8", X"FD28", X"FB25", X"FB54", X"FC4B", X"FFE2", X"00B7", X"0063", X"0200", X"01C6", X"FF26", X"0143", X"FDF3", X"FE00", X"FBB9", X"FBC0", X"F8BA", X"F8D6", X"FB1A", X"FC00", X"FCE1", X"FE29", X"0028", X"FF40", X"FD4B", X"FBA4", X"FD87", X"FC9D", X"FC19", X"FBF1", X"FAE6", X"F8D8", X"FBD8", X"FF26", X"005F", X"0209", X"0206", X"00C1", X"00CB", X"FE9D", X"FACB", X"F959", X"F97A", X"F7BC", X"F4DC", X"FA10", X"FC29", X"FB28", X"FFF3", X"FE6D", X"0097", X"006C", X"FBA3", X"F86E", X"FABE", X"F90F", X"F84D", X"FB64", X"FD87", X"FCC0", X"FD70", X"FD9B", X"FF42", X"FF80", X"FFBC", X"0063", X"FF3A", X"FD35", X"FA4B", X"F8D2", X"F8B3", X"F679", X"F663", X"F89A", X"FCB8", X"FA6A", X"FEC6", X"FFE5", X"0052", X"00C6", X"FDAA", X"FB6E", X"F974", X"F862", X"FB54", X"FBCB", X"FFC3", X"FEDE", X"FDB8", X"FC6F", X"FAAD", X"FA64", X"FA86", X"FB0B", X"FB8F", X"FA7F", X"F8D3", X"F85B", X"F812", X"F832", X"F8BD", X"FA8E", X"FD84", X"FB33", X"FF2A", X"0122", X"004F", X"FF45", X"FCAA", X"FA61", X"FD4D", X"FE55", X"0136", X"0260", X"FECA", X"FCF4", X"FC20", X"FB9C", X"F983", X"FAD8", X"F99A", X"F85C", X"F791", X"F94F", X"FB5E", X"FAF2", X"FA64", X"FADE", X"FC0D", X"FB46", X"FC9E", X"FA1C", X"FC3B", X"0005", X"0120", X"0114", X"FF59", X"FF17", X"0226", X"0683", X"0698", X"06AC", X"032F", X"FFD7", X"0153", X"FF4E", X"FEC5", X"FC2C", X"FC1D", X"FB00", X"FE10", X"FE0F", X"FDD1", X"FF03", X"005B", X"0111", X"01C1", X"FEB3", X"FC3F", X"00EE", X"FE06", X"FFAD", X"00A8", X"000E", X"FDBB", X"FEA8", X"0331", X"0897", X"05E3", X"0752", X"0381", X"034E", X"02C4", X"0427", X"02E6", X"0117", X"0125", X"0037", X"FE5C", X"FDCC", X"00BC", X"FFB0", X"02B3", X"0264", X"0230", X"0134", X"FDCD", X"00B6", X"FFFA", X"0062", X"FF4A", X"0031", X"001B", X"00FF", X"0249", X"0583", X"06F2", X"0933", X"0767", X"0772", X"04B7", X"0385", X"0039", X"01BC", X"0382", X"048E", X"013D", X"FFAB", X"0156", X"FF5F", X"FFE0", X"00BF", X"0057", X"0034", X"FEA1", X"FFED", X"00F8", X"FFBE", X"FF02", X"FF9D", X"00B3", X"00A4", X"FF92", X"0167", X"00E3", X"01D7", X"00EB", X"00ED", X"022E", X"00E3", X"FFAC", X"02F6", X"0522", X"04A8", X"0540", X"0549", X"0514", X"05F5", X"03D6", X"056E", X"02C8", X"03B9", X"0024", X"0012", X"002B", X"00A4")
--        (X"FFD3", X"FEEB", X"0073", X"0054", X"003D", X"FF8F", X"FF48", X"FE75", X"0011", X"FF8D", X"00EB", X"FDDF", X"FE63", X"FE0C", X"02D2", X"012C", X"00D1", X"FFFF", X"00B3", X"FF17", X"FFC3", X"0092", X"FE3F", X"0027", X"003B", X"0037", X"002C", X"FF03", X"FFD8", X"0016", X"FFB2", X"FFA2", X"005E", X"FF49", X"FC1E", X"FB34", X"FB04", X"FA68", X"FA26", X"F933", X"F7A7", X"F835", X"FD33", X"0183", X"0358", X"FF78", X"FBAC", X"FA30", X"FA38", X"FBFB", X"0014", X"FE36", X"0020", X"0076", X"0158", X"FF01", X"FDC8", X"FE3B", X"0060", X"0009", X"FD64", X"FBAF", X"FBB3", X"FB50", X"F8DC", X"FD18", X"FCA2", X"FBFB", X"FEAE", X"FFDD", X"FDE8", X"FEEC", X"0085", X"FFE9", X"FFB1", X"FF5D", X"FCB6", X"F91E", X"FB71", X"FBDA", X"FF6E", X"02BD", X"FFE0", X"FE76", X"015B", X"00CF", X"0153", X"0256", X"0194", X"0066", X"01AD", X"0332", X"023C", X"010F", X"0221", X"0312", X"0450", X"01A5", X"0215", X"0431", X"031B", X"01DF", X"0109", X"0102", X"FF73", X"FDE5", X"FD5F", X"FAFB", X"FD1E", X"0105", X"FE44", X"0009", X"0033", X"FFA7", X"025E", X"FF30", X"FDAB", X"03F7", X"03D8", X"037F", X"015F", X"024B", X"03BB", X"060A", X"0570", X"03F5", X"03E1", X"040C", X"02CC", X"FFCF", X"03D3", X"00DE", X"FE0C", X"FD4B", X"FBB0", X"FA9A", X"0191", X"01DE", X"FDDB", X"FD38", X"0032", X"017D", X"01B1", X"0322", X"0368", X"018C", X"015A", X"006E", X"FEB6", X"0242", X"03EC", X"03B9", X"0129", X"0108", X"0029", X"FE78", X"0249", X"0222", X"0171", X"0118", X"02A1", X"007D", X"FF25", X"FE91", X"FEC3", X"031C", X"0231", X"FE51", X"010C", X"01C6", X"FDD6", X"00A8", X"02D4", X"00BA", X"0063", X"019D", X"006C", X"02BF", X"02BE", X"0115", X"FEB3", X"012C", X"FF00", X"FF1E", X"FF68", X"0003", X"0205", X"00FA", X"0186", X"0001", X"FF6F", X"FEE3", X"0255", X"05A6", X"03E4", X"FF44", X"FE67", X"03AE", X"FE33", X"FF40", X"02CC", X"044A", X"0149", X"02AC", X"0430", X"00D5", X"0026", X"00B7", X"0153", X"FEBC", X"00CD", X"FE4D", X"FF51", X"FE07", X"FEC4", X"00DB", X"00FB", X"0031", X"01B5", X"004B", X"0330", X"0669", X"0161", X"006E", X"FEB5", X"FE45", X"FD37", X"FE5B", X"00EF", X"02E3", X"034A", X"0196", X"01C1", X"FFF2", X"FF48", X"FECF", X"FFCF", X"00DD", X"FFFF", X"FD42", X"FD9C", X"FF98", X"FF16", X"02CF", X"037D", X"02CE", X"03BA", X"027F", X"0655", X"076B", X"0545", X"029E", X"FE8F", X"FDA1", X"FF63", X"FF25", X"038D", X"00C6", X"019E", X"011B", X"0133", X"005B", X"FF58", X"016C", X"00BA", X"FFDB", X"FEFE", X"FF0C", X"FDFD", X"00A9", X"FF97", X"018B", X"024F", X"02B6", X"0330", X"049D", X"07B6", X"0C2B", X"06A0", X"01A4", X"FF75", X"FCE5", X"FF19", X"FFCA", X"0154", X"FF8C", X"00D7", X"FF22", X"FF32", X"FE11", X"FF16", X"FFF5", X"000E", X"FFF7", X"003C", X"0176", X"00B5", X"0110", X"FECA", X"0142", X"FE8D", X"FCD4", X"FC27", X"FD8B", X"050A", X"0D03", X"0793", X"0268", X"FF81", X"FCD8", X"FB5D", X"FDB4", X"FF38", X"FEEF", X"FDAB", X"FD26", X"FD44", X"FCCE", X"FD5C", X"FF57", X"025E", X"00D7", X"021A", X"017A", X"01AF", X"FF59", X"01C6", X"FE56", X"FA3F", X"F5E3", X"F39A", X"F206", X"F6D1", X"0485", X"0325", X"FFF2", X"FF62", X"FCEC", X"FA18", X"FE58", X"FCD8", X"FBA7", X"FA05", X"FC07", X"FE35", X"FD7C", X"FDB6", X"FFB3", X"012F", X"01DC", X"01F2", X"01CB", X"FDE3", X"FEDA", X"000A", X"00D4", X"FD02", X"F698", X"F30E", X"EE69", X"EBC5", X"F94E", X"FFF7", X"002F", X"0068", X"FD6A", X"FA52", X"FF76", X"FAFD", X"FA78", X"FAD7", X"FA6F", X"FD39", X"FF49", X"FF2D", X"FF7D", X"0049", X"0401", X"0341", X"FE11", X"FC4E", X"FFAC", X"00E7", X"001A", X"FC87", X"F8C5", X"F625", X"F1B3", X"EF1A", X"F7BE", X"0366", X"03A7", X"0216", X"FEA9", X"FCE7", X"011E", X"FD5B", X"FB04", X"FBBD", X"FC90", X"FDE4", X"FF88", X"FED4", X"FC71", X"FF36", X"02FA", X"0218", X"FF22", X"FF0D", X"FED9", X"FF89", X"FBB2", X"FC13", X"FC45", X"F8D8", X"F67D", X"F6A7", X"FCB8", X"0526", X"0147", X"002F", X"001F", X"018E", X"043C", X"FF8F", X"FC8C", X"FF0C", X"FB1E", X"FE21", X"FF22", X"FC4D", X"FE79", X"0111", X"0565", X"0090", X"FD8B", X"FEC0", X"FC02", X"FD3C", X"FC79", X"FC87", X"FC4A", X"F82F", X"FAC4", X"0069", X"061A", X"07F6", X"0419", X"FE35", X"01A7", X"032D", X"0812", X"0248", X"005B", X"FE26", X"F8BE", X"F91A", X"FB07", X"FA26", X"FCAD", X"FF78", X"01E7", X"FFA6", X"FDF7", X"FF16", X"029E", X"00B6", X"00F4", X"FD8D", X"00A9", X"00D1", X"0236", X"064A", X"0928", X"0A5E", X"0493", X"002E", X"00E8", X"02E3", X"0914", X"0776", X"046F", X"FF30", X"FC4B", X"F9D3", X"F83D", X"F6B5", X"F72A", X"F9FF", X"FD7E", X"FFA7", X"0087", X"00CB", X"0423", X"0397", X"05A1", X"030D", X"0494", X"040A", X"0652", X"0673", X"0761", X"092C", X"015F", X"FC3A", X"00BE", X"0247", X"09A4", X"0762", X"058E", X"0394", X"005E", X"FE27", X"FA4A", X"FA49", X"F888", X"FA2B", X"FCFA", X"0210", X"0298", X"0476", X"05CA", X"0266", X"0590", X"045B", X"02C0", X"0530", X"0823", X"0952", X"0522", X"018E", X"0344", X"FF60", X"FBC2", X"00DE", X"0764", X"07FF", X"02AB", X"0200", X"FFD4", X"0235", X"022E", X"00E2", X"FD78", X"FCCF", X"0128", X"FFDE", X"03F6", X"052E", X"0628", X"069F", X"053D", X"03EF", X"0319", X"03FB", X"07A0", X"08AA", X"076E", X"03EC", X"01B4", X"FF06", X"FCE6", X"028E", X"06D8", X"058F", X"03BD", X"044F", X"02D4", X"034F", X"031E", X"0008", X"FF51", X"FCAC", X"FD3B", X"FE48", X"00C1", X"03B7", X"06D0", X"0633", X"04C2", X"0297", X"03B1", X"06D2", X"0A16", X"07B0", X"0755", X"0136", X"0220", X"FFEA", X"00A7", X"0417", X"052D", X"0446", X"03E7", X"0261", X"009D", X"FFC5", X"0162", X"FFF3", X"FE90", X"FC66", X"FC3F", X"FE31", X"FD73", X"0150", X"038F", X"05FC", X"05FD", X"0481", X"0561", X"06A8", X"0809", X"05C5", X"064B", X"0109", X"FFDC", X"01C9", X"FFFD", X"03E3", X"05A5", X"05E2", X"0145", X"FF2B", X"006D", X"FF57", X"FFA5", X"FFBE", X"FF4F", X"FC61", X"FC33", X"FAB6", X"FB16", X"FEA1", X"026C", X"065F", X"0808", X"07BD", X"083A", X"0728", X"047F", X"04B6", X"03BA", X"01B7", X"FF6A", X"FF35", X"0033", X"02E8", X"07F1", X"059F", X"02D8", X"0163", X"011D", X"01AD", X"020F", X"013F", X"008D", X"FE3D", X"FC98", X"FBD1", X"FC8D", X"FD81", X"0227", X"05D2", X"0A82", X"0832", X"061D", X"03D7", X"0531", X"02A6", X"036D", X"0334", X"FF8F", X"FFCE", X"FEB4", X"FEE0", X"0304", X"018E", X"FDBD", X"0138", X"0270", X"023E", X"02F5", X"02A5", X"00AE", X"0190", X"01F1", X"0028", X"FC45", X"FF16", X"0175", X"06EF", X"06D6", X"059A", X"0368", X"018C", X"02EE", X"05A0", X"0320", X"026C", X"FFA1", X"0003", X"FF1C", X"0223", X"FE63", X"FCB3", X"FE72", X"00A8", X"02FB", X"03FB", X"05B2", X"0416", X"04E8", X"064B", X"0340", X"017C", X"FECC", X"FFFD", X"FFAF", X"0320", X"0312", X"003E", X"FF74", X"034C", X"01CD", X"0354", X"000E", X"02A5", X"FF71", X"FF7F", X"FFEA", X"004D", X"FF6F", X"FDF9", X"FD12", X"FBC6", X"FDBE", X"FC9D", X"FDAB", X"FC24", X"FCB6", X"FC14", X"FE09", X"FBBB", X"FDD2", X"FB5E", X"FC4C", X"FDCE", X"FE2D", X"FFBC", X"0126", X"FF2D", X"FCEA", X"FD7F", X"FF73", X"000F", X"0084", X"FEEE", X"01A9", X"0051", X"FFB6", X"0061", X"FF83", X"FE42", X"FE6C", X"FD6A", X"FE02", X"FCEF", X"FFC0", X"009A", X"FF91", X"FCA6", X"FE00", X"FCE6", X"F89A", X"F824", X"F91C", X"FB55", X"F9F9", X"FD6E", X"FC28", X"0004", X"FF3A", X"0087", X"00D3"),
--        (X"FF20", X"FF57", X"FFA0", X"00F0", X"0087", X"0181", X"00B7", X"0042", X"000B", X"FFB9", X"007C", X"0058", X"01D1", X"02AC", X"FFFF", X"FF79", X"0202", X"FF24", X"00E4", X"0077", X"0103", X"FEFA", X"00B2", X"0109", X"00DD", X"012C", X"FF00", X"FF7A", X"0005", X"002C", X"FF81", X"0182", X"FF55", X"FF89", X"028C", X"043B", X"0441", X"04CF", X"0465", X"04C6", X"0432", X"024D", X"00E6", X"04E7", X"03F8", X"0380", X"0385", X"056C", X"0473", X"0473", X"036E", X"0280", X"004B", X"FF61", X"FE93", X"01C6", X"FFD3", X"FE98", X"0169", X"FF72", X"FF59", X"00C9", X"0321", X"0795", X"0929", X"0AD8", X"0AD2", X"09B6", X"0C6C", X"07CF", X"05C5", X"05E7", X"0508", X"029B", X"044C", X"01E2", X"0522", X"0560", X"04A7", X"044F", X"02E9", X"01C4", X"00B7", X"FEA5", X"0109", X"FF7A", X"0091", X"025A", X"003D", X"FCDA", X"00BE", X"025A", X"022C", X"03DF", X"03C2", X"FF6D", X"0027", X"0180", X"FEB2", X"FFED", X"FF7B", X"FEA3", X"FE48", X"FF4D", X"FFF2", X"03B1", X"037C", X"0433", X"0405", X"007A", X"FF13", X"00A4", X"004B", X"FFFF", X"FFC2", X"FEA3", X"FDC9", X"FEFC", X"FF73", X"FEA7", X"FF5F", X"009B", X"FF59", X"FD50", X"FF57", X"FDC8", X"FF69", X"FF19", X"FF07", X"FF91", X"FF99", X"01F9", X"03AB", X"03E0", X"040F", X"052E", X"0075", X"FFC6", X"FEB0", X"0261", X"00A8", X"0124", X"0350", X"FED1", X"FFB5", X"FEAB", X"FF03", X"FD8E", X"FD28", X"FE01", X"FF9A", X"FF93", X"FE21", X"0193", X"0270", X"01EB", X"0295", X"0133", X"0252", X"046A", X"04F7", X"0575", X"04FA", X"0431", X"0321", X"FE6F", X"0292", X"022C", X"FF08", X"FF9C", X"FCBB", X"FE0D", X"FE3B", X"FB3E", X"FBF3", X"FE7D", X"FDDC", X"FC10", X"FDE9", X"FFAB", X"FE32", X"FF8D", X"FFC3", X"0060", X"FF69", X"FE90", X"00D7", X"009E", X"00D5", X"00E5", X"008C", X"FF65", X"FFE3", X"FEF0", X"0133", X"00BD", X"0100", X"002E", X"FEDA", X"F9B5", X"FAD6", X"FB4B", X"FC6D", X"FE0A", X"FD63", X"FED4", X"FFB6", X"00AF", X"0092", X"FFA1", X"FFA1", X"FDC4", X"FE86", X"FFB8", X"FE26", X"FD02", X"FE39", X"FCEE", X"FD30", X"FA0F", X"F980", X"FA59", X"FF41", X"002A", X"FD75", X"01F9", X"FF1D", X"FA28", X"FA66", X"FCD1", X"FE13", X"FE79", X"FE10", X"FFC9", X"038B", X"02C9", X"0281", X"01AA", X"FEF8", X"FF62", X"FC1B", X"FB5C", X"F910", X"FA40", X"F9DC", X"FA10", X"F96D", X"F7BE", X"F3D8", X"F4F5", X"FA1F", X"FCDE", X"FFE0", X"FEC9", X"0037", X"0032", X"FCDD", X"FE49", X"FE57", X"FD12", X"FE94", X"0112", X"010D", X"01F8", X"01EF", X"0349", X"01FE", X"FE6E", X"FB46", X"F8D4", X"F72D", X"F63E", X"F883", X"F829", X"F6B4", X"F59D", X"F486", X"F572", X"F991", X"0033", X"FEF1", X"0086", X"00DC", X"FE82", X"FA7D", X"FE21", X"FF1C", X"FEE9", X"FF89", X"FD57", X"0192", X"011B", X"FF09", X"FF0A", X"FF22", X"FC3C", X"FB5E", X"F982", X"F894", X"F938", X"F826", X"FA94", X"F948", X"FA19", X"F911", X"FBF8", X"FBFE", X"FCFC", X"00A5", X"FF9B", X"FE75", X"FBB7", X"FDA1", X"FD45", X"FBEF", X"FBF2", X"FC21", X"FB2C", X"FD78", X"FC6B", X"FA2C", X"FB81", X"FBF3", X"FA68", X"FB5D", X"F9C8", X"FB1F", X"FC0D", X"FB5F", X"FEB3", X"FE84", X"01FF", X"FFB2", X"0062", X"FA1B", X"FE8E", X"01B5", X"FFD9", X"00DB", X"F9F7", X"FCE4", X"FCCF", X"F938", X"F826", X"FB2F", X"FA00", X"F912", X"F9EF", X"FA88", X"F99D", X"FEBD", X"FE02", X"FDEE", X"FC7B", X"FCE5", X"FCFD", X"FF0B", X"01F9", X"0178", X"02C1", X"0385", X"03CF", X"FDDF", X"0439", X"FF54", X"003E", X"FFAB", X"FD5F", X"FA66", X"F977", X"F7A4", X"F88E", X"FA5E", X"F8CD", X"FC82", X"FB93", X"FD5A", X"0132", X"0131", X"0125", X"FFF3", X"FECC", X"FD1E", X"FEE3", X"FF01", X"000F", X"0168", X"032F", X"0341", X"0331", X"04A0", X"0294", X"0157", X"FEA2", X"FE05", X"FEEB", X"F909", X"FAC2", X"FBE2", X"FB4D", X"FDA9", X"FDC1", X"FEE0", X"FF34", X"FE82", X"031B", X"0547", X"0366", X"001C", X"FCB3", X"FD10", X"FF8A", X"FEE8", X"002D", X"021D", X"036B", X"0248", X"0211", X"05EA", X"02D7", X"00CA", X"FD7B", X"FD9A", X"0087", X"FAA2", X"FD66", X"00E2", X"006F", X"002C", X"FFE8", X"0025", X"00DA", X"03A8", X"04FA", X"06DC", X"032C", X"0185", X"FBB5", X"FF2F", X"FE65", X"FE93", X"0133", X"FF9C", X"00C0", X"04B5", X"05EF", X"01CA", X"0461", X"FE66", X"FD76", X"FCCB", X"01F3", X"FCE0", X"012E", X"0287", X"0153", X"FF1B", X"0224", X"051A", X"04B7", X"03F9", X"03DA", X"0607", X"0478", X"FF66", X"FD63", X"FDE2", X"FDCE", X"008A", X"009C", X"0043", X"0136", X"0371", X"07BB", X"0469", X"0455", X"FF3A", X"FE15", X"FF93", X"023C", X"FD9A", X"015D", X"03C8", X"0086", X"0172", X"02A1", X"04FE", X"04BF", X"0266", X"01FB", X"0504", X"0391", X"FD35", X"FD34", X"FE2E", X"FF5B", X"0141", X"00A6", X"00C9", X"0190", X"0397", X"083C", X"0442", X"005D", X"0041", X"FF82", X"FCEA", X"0044", X"00A4", X"FFD7", X"00CC", X"0183", X"02E7", X"0242", X"0232", X"0145", X"032D", X"03A8", X"0311", X"01CC", X"FE2A", X"FF22", X"FF93", X"FE76", X"004E", X"0051", X"0070", X"02E0", X"04BA", X"0B44", X"035D", X"030C", X"009C", X"FF49", X"0041", X"FF01", X"FEDF", X"FDFB", X"FE94", X"01DB", X"016A", X"0380", X"01ED", X"03B5", X"0159", X"029D", X"032B", X"01D2", X"FFCC", X"0102", X"FF34", X"0096", X"012B", X"FFA9", X"004A", X"0259", X"03A9", X"07CD", X"04E9", X"0352", X"010C", X"FEE8", X"FFE2", X"FEDD", X"00FE", X"FF10", X"0098", X"026E", X"01CA", X"0551", X"03F9", X"0301", X"0264", X"0116", X"FFDC", X"00F7", X"00E2", X"FFFC", X"022F", X"01C7", X"026B", X"FFD0", X"01E2", X"02F6", X"0690", X"0581", X"0413", X"FEC8", X"FE97", X"0065", X"FB54", X"FF00", X"01AE", X"FF9E", X"0088", X"028B", X"02BE", X"05A3", X"0420", X"0437", X"0512", X"0270", X"0110", X"0225", X"FF3F", X"0319", X"0554", X"02EB", X"01FD", X"0370", X"0378", X"04B7", X"0642", X"065C", X"018C", X"0029", X"FF0B", X"FF79", X"FC61", X"00FE", X"02B3", X"029F", X"0102", X"FE3A", X"0255", X"0329", X"01E2", X"0151", X"0058", X"FE56", X"FF16", X"FF47", X"0112", X"0015", X"0261", X"0335", X"0566", X"0477", X"022D", X"01E9", X"02CB", X"0507", X"02CB", X"00B6", X"FEF8", X"FFC4", X"FEE1", X"FB32", X"FFD5", X"01B3", X"FFE6", X"FD2B", X"FE2D", X"FF7C", X"FDF0", X"FE0D", X"009F", X"FF2D", X"FDDB", X"FF17", X"FF7F", X"FD46", X"FF6D", X"028A", X"013F", X"00FE", X"01AE", X"FECD", X"FECC", X"01F9", X"0387", X"0043", X"009A", X"00EB", X"00F5", X"F753", X"F9FE", X"FD47", X"FCDB", X"FA5A", X"FA52", X"F8D3", X"FA94", X"F942", X"F8E6", X"F883", X"F9A3", X"FA8A", X"F928", X"FB7B", X"FCDE", X"FBED", X"FCC2", X"FF09", X"FD65", X"FBE7", X"0156", X"0424", X"01BA", X"0074", X"FF2D", X"FF8E", X"FF6B", X"FDE6", X"FB4A", X"F9D8", X"F8F2", X"F820", X"F818", X"F83F", X"F787", X"F7BB", X"F74B", X"F560", X"F516", X"F37A", X"F43A", X"F4D9", X"F56D", X"F638", X"FA05", X"FD0A", X"FBEC", X"FB10", X"FCA5", X"0197", X"0127", X"0096", X"0085", X"0137", X"00C5", X"FEA9", X"FE8C", X"FCA9", X"FEB9", X"0053", X"FE64", X"FE7A", X"FD40", X"FA7B", X"F9A4", X"F9A4", X"F9DA", X"FA19", X"F8DF", X"F8AF", X"FA1C", X"FA42", X"FB5D", X"FB1A", X"FBE0", X"FF9A", X"013D", X"FDBB", X"FFDC", X"0062", X"FF54", X"0087", X"FF09", X"FE3C", X"FFBF", X"00B1", X"00C5", X"FFBE", X"FF9E", X"00D0", X"FF03", X"0142", X"FF8B", X"FFCC", X"FF46", X"0138", X"00CF", X"01A5", X"FE2C", X"FFD5", X"FE48", X"00C9", X"FDD8", X"0105", X"006C", X"FF43", X"0067", X"0057"),
--        (X"00C9", X"0038", X"004B", X"FF81", X"0047", X"00EA", X"FF71", X"FF60", X"FF60", X"FFAD", X"FFC7", X"0126", X"FE33", X"FFB5", X"01BC", X"FFD3", X"FF1A", X"0004", X"0128", X"FFCA", X"FE7C", X"FF5F", X"0060", X"FE7B", X"0024", X"006F", X"00FD", X"0219", X"022B", X"007E", X"0184", X"FF0A", X"FFD7", X"FEE9", X"FCC8", X"FE1C", X"FD6A", X"FE65", X"FDC1", X"FD66", X"FC4F", X"FDA9", X"FEEC", X"FCE8", X"FC4D", X"FB80", X"F984", X"FB7A", X"FAF9", X"FCED", X"FDE3", X"FE1C", X"00E5", X"0038", X"FF9D", X"FF7C", X"FE77", X"FF1A", X"FFB5", X"FFB4", X"FDB9", X"FCE4", X"FCC3", X"FC5E", X"FC0A", X"FE44", X"FBF6", X"FBDC", X"FE0F", X"FDF9", X"FDAA", X"FD04", X"FDB0", X"FE8E", X"FB6D", X"F9FD", X"FA3C", X"F872", X"FAD1", X"FA9B", X"FED7", X"0046", X"0020", X"00F3", X"FED2", X"0137", X"0031", X"FC0C", X"006C", X"FB20", X"FC3D", X"FF58", X"FD2E", X"FAD2", X"FC8E", X"FC27", X"FA5C", X"FA55", X"FB03", X"F8A3", X"FAE0", X"FB45", X"FD0D", X"F9D7", X"F9D2", X"FC13", X"FC37", X"0017", X"000D", X"0235", X"01E1", X"FFD4", X"014B", X"FFA4", X"FE67", X"FCD9", X"FE14", X"003C", X"0081", X"015C", X"FF5A", X"FDFA", X"FDA7", X"FFC9", X"FE95", X"FD45", X"FDD7", X"FEDE", X"FCFA", X"FDD4", X"FC1B", X"FB2D", X"FC9F", X"FFD4", X"00E2", X"01D4", X"041D", X"03E8", X"FF95", X"001B", X"FE46", X"FEFD", X"FED0", X"03F3", X"FEBF", X"0134", X"01D5", X"01AD", X"0072", X"00DD", X"009B", X"067B", X"041F", X"0328", X"03EF", X"0603", X"03F9", X"053D", X"03A5", X"05E3", X"05FE", X"05BB", X"0835", X"0971", X"0772", X"04E0", X"013C", X"FFAF", X"FFB7", X"0086", X"FEAA", X"FD01", X"FC7B", X"FE5C", X"FF01", X"FED4", X"FE8F", X"FDB7", X"FFFB", X"0034", X"0010", X"020A", X"00A8", X"0221", X"033E", X"023B", X"05EB", X"0514", X"074D", X"0528", X"080B", X"094F", X"09B7", X"086E", X"04B6", X"02E6", X"0010", X"FDCC", X"FC2C", X"FB54", X"FDA0", X"FEF9", X"FE5C", X"FD49", X"FE61", X"FE55", X"FCE9", X"FE9F", X"FEFA", X"FF60", X"FF83", X"0068", X"02FA", X"0209", X"0494", X"04B5", X"04EA", X"0462", X"05FA", X"0722", X"0878", X"08FA", X"05E1", X"033C", X"026C", X"FBF4", X"FB7C", X"FBA2", X"FDA4", X"FF42", X"FE02", X"FCAB", X"FD39", X"FE48", X"FC38", X"FD8A", X"FC3A", X"FD71", X"FC71", X"FDF1", X"0068", X"03A0", X"0686", X"04CB", X"0428", X"041F", X"027C", X"02F0", X"0721", X"0A2E", X"0599", X"0224", X"006F", X"FEB3", X"FEA7", X"FCE9", X"FB0C", X"FC43", X"FDF8", X"FD5C", X"FE3A", X"FCF8", X"FE15", X"FD38", X"FDC4", X"FDE3", X"FA7B", X"FDE4", X"0069", X"0415", X"048A", X"03E3", X"02E4", X"00BA", X"0251", X"036D", X"0347", X"0614", X"02DE", X"FE63", X"002A", X"FCD7", X"F8C3", X"FD2D", X"FE2A", X"FD36", X"FEA0", X"FE2F", X"FE2D", X"FF43", X"FE43", X"FF4A", X"FFC8", X"F9DE", X"F81E", X"FB2E", X"0028", X"00D5", X"02D8", X"0297", X"FF5C", X"FFF4", X"FF9E", X"0034", X"01BC", X"036C", X"01EA", X"001E", X"FEFD", X"FC76", X"FA07", X"FAEA", X"FB31", X"FE88", X"FE97", X"FCE9", X"FF99", X"FF25", X"FF48", X"FECF", X"FD09", X"FA40", X"F88C", X"FDAA", X"FE72", X"0011", X"FF2C", X"00E5", X"FF96", X"FEE3", X"FED7", X"FBCF", X"FEC4", X"03C7", X"0624", X"0159", X"FF0B", X"FC77", X"F830", X"FBE3", X"FC1B", X"FDF8", X"FF57", X"FBE4", X"FD49", X"FFD2", X"FF79", X"0066", X"015B", X"0298", X"0222", X"FFD4", X"FCFE", X"FC76", X"FD52", X"002E", X"01CF", X"FE69", X"FC8A", X"FCC9", X"FC51", X"FF6D", X"03D5", X"FD71", X"FFCD", X"FF68", X"FB12", X"FCAE", X"FC88", X"FDB1", X"FEFE", X"0009", X"FFDB", X"01D9", X"0189", X"047C", X"06F6", X"0719", X"0485", X"019F", X"FE8D", X"FE3E", X"FF7A", X"00CB", X"002D", X"FEA4", X"FAB8", X"F82E", X"FB89", X"0117", X"04B7", X"0500", X"FF55", X"FDEC", X"FAE3", X"FCB4", X"FEAE", X"FE33", X"FF96", X"00D9", X"00F8", X"037B", X"042E", X"051E", X"06DB", X"065E", X"02F1", X"01CD", X"FF8D", X"00B6", X"FF1C", X"FE35", X"FC65", X"FBC2", X"FA69", X"FA8E", X"FC85", X"00A4", X"056C", X"02ED", X"FFA8", X"FF8D", X"FC9E", X"0006", X"0253", X"009C", X"FFC0", X"0253", X"04BA", X"05CE", X"03AF", X"02BC", X"0608", X"0301", X"00D6", X"0075", X"03BC", X"FF75", X"FDCB", X"FB60", X"FC8E", X"FB76", X"FE08", X"FF77", X"FFCF", X"FFB5", X"08D3", X"03FC", X"FF19", X"FFF9", X"FC4F", X"00E2", X"03F9", X"017F", X"0058", X"01E4", X"0577", X"042E", X"04B9", X"034E", X"03CC", X"0284", X"FF04", X"014C", X"03AC", X"02F6", X"FDA8", X"FD44", X"FB94", X"FDF1", X"0007", X"FF2F", X"0098", X"01D3", X"078F", X"0062", X"FF2C", X"FF26", X"FD50", X"03E9", X"056C", X"0267", X"0142", X"0478", X"054B", X"0575", X"02ED", X"01A3", X"02F6", X"FF92", X"FF70", X"00EE", X"025B", X"0162", X"0006", X"0054", X"FE4C", X"FEF1", X"FD2E", X"FE62", X"FE14", X"FD97", X"039B", X"01C1", X"FC94", X"FF69", X"FD13", X"030A", X"0305", X"05A8", X"04E0", X"0452", X"0517", X"0436", X"03D9", X"0250", X"FE7A", X"FD02", X"FD3E", X"00A0", X"00F2", X"FFC6", X"FEDE", X"002F", X"0118", X"FDCA", X"FE5E", X"FE49", X"FE67", X"FE46", X"0107", X"0121", X"014E", X"FC1E", X"FD59", X"04C9", X"02F4", X"062B", X"05AC", X"0475", X"04FD", X"024C", X"0040", X"FE5E", X"FA40", X"FA75", X"F9FF", X"FD5D", X"FD61", X"FDAC", X"FE2E", X"FEA4", X"FF60", X"0091", X"011A", X"0184", X"FFFC", X"011C", X"0351", X"034E", X"FFDD", X"0322", X"0101", X"047C", X"05D0", X"05D5", X"0462", X"04FE", X"03B3", X"0152", X"FE12", X"FBFB", X"FA6D", X"F9C0", X"FADF", X"FBD1", X"FEF7", X"FF94", X"FFB8", X"0085", X"03E7", X"03CC", X"045D", X"02ED", X"0381", X"02F3", X"FE53", X"FEB2", X"FF0C", X"FF94", X"034A", X"019B", X"056B", X"07C5", X"05E1", X"059A", X"0348", X"01B9", X"FD0E", X"F96A", X"FA39", X"F946", X"FB8B", X"FB89", X"FCC4", X"FDEE", X"0114", X"0352", X"06A5", X"0517", X"06EE", X"0879", X"02FF", X"00FB", X"FEF4", X"00D4", X"0056", X"FFAB", X"016D", X"0189", X"0305", X"0229", X"05DB", X"05B4", X"05F0", X"03BD", X"0110", X"0159", X"FF27", X"0065", X"017B", X"0068", X"01DD", X"036B", X"05AC", X"04AC", X"078A", X"081E", X"08A4", X"0A4A", X"0873", X"0111", X"FECE", X"FFC1", X"00DD", X"FF88", X"00E4", X"0196", X"FEBA", X"FDF1", X"FE38", X"00BD", X"06BE", X"0510", X"05CB", X"05AF", X"04E4", X"053C", X"040A", X"0462", X"05E5", X"0434", X"08F8", X"06BF", X"0854", X"0964", X"08A6", X"0B4E", X"05CA", X"0368", X"FEF0", X"006D", X"FFB1", X"000E", X"FD75", X"FC69", X"FB1E", X"F8E9", X"FA10", X"FB39", X"FE58", X"FFFB", X"0062", X"01D0", X"021F", X"0182", X"0259", X"023A", X"0445", X"0445", X"056D", X"05CC", X"07E9", X"08E1", X"0804", X"09D4", X"05B7", X"0172", X"FDF6", X"FF61", X"FEDB", X"017B", X"01B5", X"FDCD", X"FD99", X"FCDD", X"FC73", X"FA95", X"F950", X"FC2F", X"FE94", X"FBDB", X"FA1B", X"FC77", X"FD6F", X"FB58", X"FC9A", X"FF20", X"FF92", X"00BB", X"0301", X"04E6", X"04B2", X"0414", X"FEA2", X"0180", X"006C", X"0180", X"00C7", X"FEF7", X"004D", X"01CF", X"0281", X"FEDF", X"007A", X"0008", X"FDE0", X"0012", X"FFC2", X"FE15", X"FF5F", X"FDB0", X"FE3B", X"FB91", X"FD31", X"FBE4", X"F923", X"F9AD", X"FFB8", X"0104", X"FD57", X"0052", X"0035", X"FE3E", X"FFEF", X"FF5B", X"FF86", X"FEF1", X"003A", X"FEC6", X"0034", X"FF1D", X"0048", X"FF6F", X"FEC3", X"FFA5", X"FF63", X"FE97", X"0035", X"FBD0", X"FD73", X"FD1F", X"FCDB", X"FE84", X"FD02", X"FC8B", X"FEB6", X"FC78", X"FDAA", X"FC4F", X"FEE8", X"0038", X"005D", X"00E9"),
--        (X"FF9B", X"FFB3", X"00A7", X"FEC7", X"000B", X"FFF7", X"0099", X"014F", X"FE23", X"0029", X"0014", X"FEA7", X"FE63", X"FF83", X"FFE0", X"0012", X"FF0E", X"0102", X"FFAB", X"FF29", X"FEC3", X"FFEF", X"FFE5", X"0049", X"FFF2", X"FFF8", X"FF38", X"FE19", X"00AA", X"00A9", X"0069", X"0095", X"0063", X"007D", X"0237", X"FFC5", X"FC73", X"FCE2", X"FDD9", X"FCD0", X"FDFA", X"FBB2", X"FE9F", X"0158", X"007F", X"FD3E", X"FCAB", X"FE92", X"FF82", X"00F4", X"00F5", X"00FC", X"0050", X"FF9D", X"FFC9", X"00A0", X"0010", X"FFEB", X"FEA0", X"FF3B", X"FFB4", X"FF7E", X"FDAA", X"FE06", X"FE33", X"FEE2", X"FC1D", X"FA5B", X"F9EC", X"F8E5", X"F816", X"FB3A", X"FD85", X"FDF5", X"0068", X"FED3", X"FE0F", X"FDE3", X"FCD9", X"FDDA", X"FE79", X"0096", X"01A1", X"0050", X"FF6B", X"FF9F", X"FFEC", X"018A", X"FFBA", X"FF61", X"FFF3", X"00EB", X"01D3", X"0233", X"010E", X"FF16", X"01D7", X"FF34", X"FE8E", X"0252", X"0081", X"00B3", X"016F", X"008F", X"FFC7", X"FED4", X"FED0", X"FE98", X"FD36", X"003B", X"FEF2", X"FF07", X"001B", X"FF9B", X"FEEA", X"02B4", X"FF34", X"00D3", X"0163", X"01E9", X"01BB", X"03F9", X"051B", X"043A", X"0536", X"FF87", X"0207", X"02FE", X"FF9B", X"FE1E", X"FF39", X"FCB9", X"FBFD", X"FCBC", X"FC9A", X"FDF6", X"0126", X"0134", X"01DC", X"FF6E", X"00A1", X"FF73", X"FED2", X"00B8", X"FCFA", X"FED6", X"FC02", X"FCC9", X"FD36", X"FED9", X"0203", X"054E", X"0546", X"073F", X"03E2", X"021A", X"FF62", X"FF8D", X"FD85", X"FD9D", X"FE81", X"FF1D", X"0015", X"FD2B", X"FEC4", X"0132", X"006C", X"FFCF", X"FF37", X"FFCE", X"FD0E", X"FD10", X"F9C8", X"F68F", X"F72A", X"FA6A", X"FBAC", X"FFDF", X"0387", X"05B6", X"0532", X"04E6", X"073D", X"0889", X"06B3", X"03C5", X"0693", X"02FB", X"035C", X"FEFE", X"FE4E", X"FD34", X"005C", X"0386", X"0100", X"0005", X"0041", X"FD23", X"FA28", X"F8AA", X"F4BD", X"F5F1", X"F9ED", X"F9F9", X"FED0", X"FEEC", X"02F6", X"0436", X"02B9", X"06B0", X"072A", X"07A0", X"085F", X"04D2", X"0350", X"0344", X"0349", X"003F", X"FD59", X"FD50", X"01F5", X"0518", X"0268", X"00E9", X"FD17", X"FB34", X"F86F", X"F890", X"F8D2", X"F964", X"FBEF", X"FD50", X"FF7D", X"FEA9", X"0003", X"0193", X"0233", X"04C7", X"08F3", X"04E4", X"02A6", X"017A", X"0134", X"00FB", X"FFC2", X"00C8", X"FF0E", X"0002", X"041C", X"06B8", X"048F", X"0377", X"FF21", X"FC4F", X"FA57", X"FB0C", X"F93F", X"FD4C", X"00B1", X"FFB7", X"FF1B", X"FFBE", X"FF16", X"FFE4", X"FF54", X"0178", X"058D", X"032F", X"FCA2", X"FC63", X"FD05", X"FE79", X"FE48", X"FF9A", X"FE33", X"00FF", X"07D9", X"09F4", X"0801", X"02F4", X"FFE4", X"FC94", X"F8B1", X"FCCA", X"FE55", X"0186", X"024D", X"00F9", X"FF76", X"FF30", X"FEB0", X"FED5", X"FDD2", X"FF39", X"041D", X"0194", X"FB87", X"FCC4", X"FEA0", X"FD92", X"FD59", X"FEC2", X"FD21", X"01F1", X"075E", X"0DCC", X"09D6", X"03D5", X"FF3B", X"FA2D", X"F796", X"FB94", X"005D", X"0470", X"02BF", X"01F7", X"0071", X"FD7B", X"FC5F", X"FC7D", X"FA52", X"01ED", X"0A11", X"0459", X"FED2", X"FDA3", X"FF17", X"FF0A", X"FFDA", X"FE1D", X"FE1C", X"FFDE", X"069C", X"0C03", X"086C", X"0221", X"FEC7", X"FAC9", X"F8EC", X"FF53", X"0625", X"0694", X"0143", X"010E", X"FCC3", X"FD9A", X"FB4D", X"FA28", X"F786", X"02EA", X"09FE", X"05E3", X"FE4F", X"FEDA", X"00A4", X"01DC", X"01F8", X"FF4B", X"FC7D", X"FB9E", X"FCCF", X"041E", X"06DD", X"01A7", X"FFAF", X"FCFF", X"FA71", X"00C1", X"04F0", X"0239", X"FDFC", X"FD7E", X"FF38", X"FC39", X"FB31", X"F8B6", X"FDC3", X"070E", X"0928", X"03B6", X"00DF", X"FE99", X"0115", X"0281", X"01B3", X"FF95", X"FCBB", X"F809", X"F858", X"FDE6", X"0467", X"03E7", X"016E", X"FE40", X"FBD6", X"01C7", X"FFF4", X"FD0D", X"FD0C", X"FED1", X"FCEE", X"FC58", X"FB6B", X"F9E7", X"FFF5", X"0695", X"06D3", X"031B", X"FEA3", X"FD4D", X"FFA1", X"FFB2", X"009A", X"FE29", X"FB32", X"F9C0", X"FA92", X"FDEC", X"05BB", X"0108", X"0110", X"00C3", X"FD25", X"FE0B", X"FDDC", X"FA43", X"FE16", X"FD19", X"FDD4", X"FBB6", X"FC93", X"FDB8", X"0533", X"06E7", X"03BA", X"0037", X"FDB7", X"FD72", X"FFC1", X"FE78", X"FF95", X"FC96", X"F929", X"F956", X"FD95", X"FE2A", X"00BE", X"021B", X"FFE8", X"001A", X"FE81", X"FFA7", X"00C2", X"FD8B", X"FE48", X"FD4A", X"FC89", X"FCE9", X"FF7F", X"024E", X"069E", X"070B", X"00CA", X"FBC2", X"FBE3", X"FC94", X"FC64", X"FD0F", X"FB8D", X"FA8E", X"FAE2", X"FCE3", X"FFFA", X"FE3A", X"FF3C", X"0113", X"FEC2", X"FFBC", X"FCB0", X"0222", X"0035", X"FCD6", X"0019", X"FDFB", X"FC1B", X"FE3F", X"001E", X"0506", X"08F2", X"042D", X"FF53", X"FC76", X"FD7B", X"FCE3", X"FD01", X"FF83", X"FC1B", X"F9EA", X"FA96", X"FF8A", X"01D8", X"FF64", X"013F", X"00C9", X"004A", X"015E", X"FEAA", X"01A5", X"FE35", X"FFA8", X"0363", X"FF24", X"FC50", X"FF47", X"032A", X"05D5", X"05EC", X"029D", X"FFBF", X"FE5E", X"FF1B", X"FEB6", X"FD29", X"FE68", X"FD64", X"FE72", X"FF61", X"0180", X"0370", X"01B4", X"FFCC", X"012E", X"FFDE", X"FDC4", X"FFE6", X"0138", X"FF07", X"0157", X"0223", X"0047", X"0127", X"FF9D", X"02AD", X"0375", X"02E5", X"005B", X"FDEB", X"FE34", X"FE74", X"FDF1", X"FFC9", X"FFAB", X"007C", X"016C", X"05B9", X"0575", X"04DC", X"04F0", X"0169", X"00C5", X"00E2", X"FC52", X"FDFD", X"024A", X"00CC", X"01D5", X"03CF", X"008E", X"01C3", X"01E3", X"FF8F", X"FFEE", X"0052", X"FFE1", X"FD10", X"FFC7", X"006F", X"0068", X"FFD7", X"0213", X"038D", X"0228", X"0612", X"07C4", X"05AE", X"04B5", X"FE7F", X"FFE9", X"FF52", X"FF1A", X"FF4F", X"0175", X"028A", X"02C6", X"041A", X"027F", X"FFCF", X"FEF5", X"FF22", X"FC77", X"FDF2", X"FF97", X"FFCE", X"FFA4", X"003A", X"0037", X"021A", X"017C", X"01D5", X"02E5", X"0422", X"0544", X"03C1", X"0492", X"FCD1", X"FF5E", X"010D", X"FF24", X"0197", X"02AB", X"0386", X"00EA", X"01B8", X"004A", X"006B", X"007D", X"FE7E", X"FF14", X"FEF8", X"000D", X"01DB", X"FFF3", X"0128", X"00F2", X"005E", X"FEDA", X"011F", X"01AC", X"04F4", X"0708", X"0569", X"0226", X"FE07", X"FFA7", X"0126", X"016D", X"01A1", X"02D7", X"011E", X"0091", X"FC5B", X"FCB8", X"FFDB", X"FD63", X"FED5", X"FFDC", X"0065", X"01BE", X"0177", X"0149", X"0137", X"FFFF", X"FFC0", X"0044", X"0270", X"00D1", X"03E3", X"04F8", X"04FF", X"01F6", X"FDF7", X"FF86", X"0164", X"FEF5", X"FDDE", X"FDF5", X"0076", X"015A", X"FFEB", X"FFF8", X"0164", X"01F2", X"018D", X"00D4", X"031C", X"0118", X"012A", X"01BC", X"0131", X"01B1", X"0038", X"009E", X"0259", X"03F0", X"0487", X"0434", X"044C", X"FF0B", X"FEE1", X"FF2C", X"FF34", X"FED6", X"00DF", X"FECF", X"FF03", X"032C", X"02DA", X"0546", X"047B", X"02D3", X"0511", X"052A", X"070D", X"0464", X"03AC", X"033C", X"017D", X"0285", X"044A", X"0636", X"061C", X"08AD", X"04DA", X"0443", X"045B", X"01A8", X"FF06", X"FEF7", X"00B7", X"FFDE", X"FF4F", X"0200", X"019D", X"0263", X"0242", X"0372", X"028F", X"057D", X"075F", X"056E", X"068E", X"0643", X"0765", X"0459", X"0475", X"04EE", X"051B", X"02E0", X"048A", X"063C", X"034F", X"03D7", X"0260", X"FE58", X"FFC1", X"FF06", X"0028", X"FF26", X"00BF", X"00ED", X"FE6D", X"FCB9", X"FF13", X"FFA4", X"FE9B", X"FED0", X"FF9E", X"FF5A", X"020A", X"FC5A", X"01D6", X"FE3E", X"FE3E", X"FF1B", X"FF0D", X"FF69", X"FE23", X"FD17", X"006D", X"FC1B", X"0185", X"0140", X"FF2A", X"FF9D"),
--        (X"FF79", X"FF22", X"004F", X"FF2F", X"0117", X"0154", X"FF30", X"FFF6", X"FF0E", X"FF2F", X"004D", X"0027", X"0033", X"016C", X"FF46", X"00F5", X"005F", X"FF67", X"00DC", X"0055", X"FF5D", X"FEC0", X"FF4E", X"013B", X"00E5", X"FFE3", X"FFF3", X"00B4", X"00EB", X"FFC3", X"0032", X"00B0", X"008C", X"00E1", X"00C5", X"0062", X"007B", X"0081", X"012A", X"FFFE", X"FFDB", X"0120", X"0175", X"FFB9", X"0071", X"FFC3", X"001F", X"FF23", X"014A", X"0018", X"001F", X"0049", X"00AB", X"FF76", X"FF4F", X"00D7", X"00A1", X"FFC8", X"FFDF", X"FFA6", X"FE4C", X"0156", X"0283", X"02A2", X"03CD", X"0606", X"07B7", X"075E", X"045F", X"0723", X"09F8", X"0819", X"02ED", X"011E", X"FEBB", X"0098", X"FEC7", X"FE97", X"FF2A", X"FF65", X"FF73", X"FD9D", X"01B0", X"0014", X"0021", X"00C4", X"012F", X"FEBC", X"00A3", X"043E", X"03D5", X"0346", X"023B", X"0713", X"025B", X"021E", X"FF57", X"0079", X"00A4", X"0044", X"0105", X"00D5", X"00B9", X"007F", X"FD77", X"FF9F", X"FFE9", X"FDAC", X"FF1E", X"FCCF", X"FE83", X"FF60", X"00EA", X"012E", X"FF3D", X"FC8C", X"017E", X"0580", X"05C0", X"03B8", X"041D", X"0402", X"01CC", X"FFC2", X"FE9E", X"FF95", X"FE65", X"FBD7", X"FCA6", X"FEF8", X"FE9C", X"0048", X"00A8", X"00FD", X"013E", X"FF67", X"FC34", X"FAA4", X"FB36", X"0087", X"FF66", X"0056", X"0266", X"FE34", X"054A", X"0475", X"0397", X"FE00", X"FF57", X"FDF7", X"FE33", X"FC7B", X"FB30", X"FC30", X"FAA7", X"FB53", X"F977", X"FAF4", X"FF50", X"FDED", X"0052", X"FF23", X"004E", X"01C5", X"FF29", X"F9FF", X"FC87", X"0223", X"016E", X"FF5F", X"FE50", X"FCE6", X"0316", X"FC06", X"FB36", X"F9C7", X"F77B", X"F725", X"FA09", X"FB6C", X"FB9A", X"FA38", X"FD73", X"FC73", X"FC8F", X"FC00", X"FEDC", X"FDB5", X"FE20", X"FD3A", X"FF81", X"FF8D", X"FFD7", X"FB94", X"FF2E", X"FFC7", X"FE6D", X"FC89", X"FF43", X"F95D", X"FB8D", X"F8EB", X"F767", X"F5A8", X"F461", X"F7D2", X"F91B", X"FAA9", X"FC6A", X"FEC6", X"019B", X"FE8E", X"FEFB", X"FF07", X"FF63", X"FDAA", X"FF84", X"FEE0", X"FDD0", X"FDF7", X"FCDD", X"FCFF", X"00FA", X"FF23", X"0061", X"FB96", X"FCBC", X"F885", X"F8FC", X"F7AC", X"F7A0", X"F635", X"F7AD", X"F82A", X"FA62", X"FDFE", X"FE30", X"FEE9", X"01EA", X"0022", X"FCF0", X"FD7C", X"FCC4", X"FF25", X"FCF0", X"FB34", X"FC87", X"FAFF", X"FCD0", X"FDE9", X"FA05", X"FC49", X"FEDB", X"FBA2", X"FBC2", X"F8FF", X"F9D9", X"F888", X"F7FB", X"F7E5", X"F98D", X"FB3E", X"FE19", X"FF14", X"0126", X"008B", X"00CD", X"0063", X"FEDB", X"FBE3", X"FD02", X"FC8B", X"FBD9", X"FA6B", X"F9F3", X"F71C", X"F90B", X"F81C", X"F781", X"FD9D", X"FF0A", X"FC9A", X"F83C", X"F8B9", X"F808", X"FB41", X"FB49", X"FCF8", X"FE67", X"FE80", X"FF36", X"FE8D", X"FED2", X"FC12", X"FE56", X"018F", X"FDC5", X"FBDB", X"FD4B", X"FCC7", X"FB99", X"F956", X"F772", X"F7E9", X"F88C", X"F701", X"FA88", X"FF13", X"FE33", X"FCDE", X"F7D4", X"F9D2", X"FAFA", X"FE49", X"FDA5", X"FE26", X"FF17", X"FE3B", X"FE24", X"FE3C", X"FF6B", X"FBF5", X"FFFF", X"028C", X"00B5", X"FDA7", X"FE3B", X"0155", X"FF9B", X"FEC9", X"FB7F", X"FC7A", X"F98C", X"F927", X"FB84", X"0198", X"001E", X"F9B8", X"F7B8", X"F921", X"FF37", X"FF9A", X"0106", X"0008", X"00DB", X"0012", X"FF83", X"FF90", X"0060", X"0026", X"061B", X"0454", X"00F8", X"FE9A", X"0004", X"0296", X"0177", X"0333", X"01C3", X"FF8B", X"FE34", X"FC81", X"FAFE", X"0275", X"FF2B", X"FDA9", X"FA42", X"FCA6", X"00F2", X"02CD", X"0525", X"05AB", X"0314", X"015F", X"01EF", X"0263", X"03D5", X"06F3", X"082B", X"0384", X"030D", X"FFF0", X"006A", X"0306", X"00B6", X"039E", X"017B", X"0420", X"01DD", X"0055", X"FE11", X"FEF0", X"FFA0", X"FE08", X"FBD9", X"01A2", X"0437", X"0590", X"090E", X"0682", X"04D7", X"05E2", X"03D8", X"031A", X"0593", X"06BE", X"03F8", X"038E", X"037C", X"0063", X"00A8", X"0152", X"021A", X"0110", X"01ED", X"0231", X"0286", X"0281", X"FFF2", X"01F5", X"FEA9", X"FF70", X"FE2A", X"02AA", X"0164", X"0700", X"0735", X"07DF", X"069D", X"039C", X"0634", X"0566", X"044B", X"01E3", X"044A", X"03DE", X"043B", X"0047", X"0084", X"012C", X"FEF7", X"000B", X"019E", X"00CC", X"0272", X"0326", X"FD65", X"0204", X"FEE7", X"FEAF", X"FE80", X"00FA", X"FF93", X"0584", X"076E", X"079A", X"067F", X"0574", X"0552", X"03B5", X"0062", X"02FD", X"0539", X"02B7", X"036B", X"007F", X"FF6C", X"FE7A", X"FF01", X"00D0", X"0169", X"FFAF", X"025E", X"045F", X"0147", X"0176", X"007B", X"FFE5", X"FF63", X"FF05", X"FEA0", X"022F", X"031C", X"06D1", X"06E4", X"047F", X"0585", X"0239", X"029D", X"03CF", X"0651", X"0410", X"0065", X"FDCB", X"FE87", X"FEA2", X"FF56", X"01BB", X"029A", X"FEB9", X"FE6F", X"03BF", X"0159", X"FF6B", X"FD91", X"FFC8", X"FC36", X"FECB", X"FE72", X"FD66", X"FE01", X"0329", X"034D", X"0487", X"046A", X"0260", X"03D8", X"04DC", X"0614", X"03AE", X"0112", X"FEFE", X"FF83", X"0174", X"FF9A", X"02E4", X"0089", X"01EC", X"0196", X"0736", X"025F", X"04E1", X"00E8", X"FC8A", X"FC40", X"0003", X"0076", X"FAFA", X"F9F2", X"FEDE", X"003D", X"02BC", X"023F", X"02EB", X"0225", X"0413", X"02E6", X"0163", X"011F", X"FFE7", X"0019", X"0243", X"01DA", X"024B", X"0236", X"0083", X"030B", X"0602", X"02C7", X"040A", X"FE6C", X"0089", X"FCA1", X"FE9A", X"FE51", X"F97A", X"FBEB", X"FB52", X"FD7A", X"FCFF", X"FF37", X"02AC", X"00E4", X"FFFC", X"0003", X"FD91", X"019A", X"FFEE", X"0234", X"0103", X"0371", X"FEBB", X"FE16", X"FC4A", X"03D6", X"0781", X"0336", X"FFBA", X"00D1", X"0086", X"FD90", X"FF2F", X"FCBF", X"FAFA", X"F8C8", X"F9F6", X"FC99", X"FDD4", X"FC0C", X"FBF2", X"FBE5", X"FD23", X"FE1E", X"FE6D", X"FE44", X"FE21", X"00AE", X"023D", X"0048", X"FDC6", X"FB48", X"FC8A", X"04CC", X"03D2", X"02E6", X"0040", X"0195", X"010D", X"FDF7", X"FF15", X"FEF0", X"001E", X"FB24", X"F98E", X"F7BE", X"FA2C", X"FAA9", X"F7AC", X"F941", X"FA1A", X"F860", X"F9B9", X"FCF2", X"FD3B", X"FFD0", X"FEEB", X"FF74", X"FF0B", X"FD5A", X"FEC7", X"010B", X"00A2", X"FF99", X"00C0", X"005C", X"FFDA", X"FDEF", X"FD46", X"FDDE", X"013B", X"FF20", X"FCD1", X"FCE3", X"FAA2", X"F836", X"F951", X"FA0F", X"F865", X"FA77", X"FB32", X"FB73", X"FDDE", X"FF3B", X"022A", X"02D1", X"01CF", X"0019", X"FE04", X"01BD", X"00A2", X"02FD", X"FE97", X"00B7", X"FFDC", X"FE12", X"FA00", X"FD87", X"014B", X"00B6", X"FFEE", X"002E", X"FD2D", X"FCF1", X"FBA1", X"FC86", X"F9BF", X"F8FB", X"F991", X"FA6D", X"FD85", X"FE86", X"01DB", X"052A", X"0510", X"02F7", X"0215", X"FEF3", X"044D", X"0149", X"FFF9", X"0229", X"FF30", X"00EB", X"FD6C", X"FD59", X"018D", X"0025", X"FFF2", X"0328", X"FF8D", X"FFFA", X"FC0E", X"FD5C", X"FDD8", X"FF90", X"FB09", X"FD77", X"FDF0", X"FE2C", X"0068", X"0705", X"05E6", X"0050", X"FF50", X"FD37", X"00EF", X"0098", X"00EB", X"0160", X"0083", X"022A", X"020D", X"0423", X"030E", X"033C", X"0308", X"00F5", X"003B", X"0121", X"020C", X"0396", X"004D", X"0112", X"FDDD", X"FE7A", X"FD5E", X"FB63", X"FC20", X"0136", X"026D", X"FFDA", X"0099", X"0145", X"FEF3", X"00CA", X"FEED", X"00CA", X"FFD8", X"FF1D", X"0070", X"FE59", X"FDFD", X"FE36", X"FD8A", X"FC4B", X"FD1D", X"FB90", X"0013", X"FFA4", X"FACD", X"FDE2", X"FF86", X"FC05", X"FA34", X"FD2B", X"FC28", X"0062", X"FF25", X"FF7B", X"FB96", X"0153", X"00B0", X"FEEF", X"FF7C"),
--        (X"00AD", X"FF45", X"0039", X"FE78", X"002A", X"007B", X"00D7", X"0033", X"0027", X"00C0", X"00E7", X"0015", X"00D5", X"00F6", X"FF49", X"00C1", X"007A", X"FEC2", X"FFE5", X"0035", X"FFE4", X"FF5D", X"013B", X"FFB3", X"FF7B", X"FF79", X"FE84", X"FE3A", X"FF55", X"FFC1", X"00BD", X"FEEF", X"00BC", X"002C", X"FEE8", X"FF9E", X"0186", X"00F4", X"02A3", X"023C", X"0288", X"023A", X"00E6", X"FDB8", X"FFEB", X"01C9", X"FFD2", X"FFAE", X"0095", X"FED6", X"FDC3", X"FED2", X"FEC9", X"FFD7", X"FFAD", X"004A", X"FFB4", X"FEE8", X"00AF", X"0012", X"FF02", X"FFA3", X"0087", X"0151", X"03A6", X"052C", X"024C", X"037C", X"022D", X"00AC", X"0046", X"FF09", X"0031", X"04A8", X"035C", X"059F", X"02DF", X"0379", X"FEA4", X"FF0F", X"0049", X"FF27", X"FFA1", X"FF15", X"FF5D", X"FE20", X"FEAF", X"FD4C", X"00C5", X"0125", X"0009", X"0265", X"0524", X"0654", X"07A0", X"07E3", X"0375", X"034A", X"0485", X"0314", X"02A9", X"040E", X"03B3", X"065B", X"0611", X"043C", X"02A1", X"FFED", X"0165", X"0093", X"0094", X"FDA0", X"FF5F", X"00A6", X"FF1D", X"FC80", X"FFF5", X"0589", X"0408", X"04F4", X"0726", X"074E", X"047B", X"0688", X"049E", X"040D", X"04A0", X"04DF", X"081B", X"078D", X"0504", X"03D6", X"007B", X"FDF8", X"0193", X"0176", X"02E6", X"009F", X"FDD4", X"FE4E", X"FFF1", X"00D6", X"FDBB", X"0052", X"045D", X"00E4", X"0324", X"0465", X"05CD", X"062F", X"0338", X"FF01", X"FC93", X"FC53", X"FD99", X"FFA2", X"0353", X"03BB", X"0479", X"022A", X"011B", X"0254", X"02A7", X"04E4", X"03F4", X"00A0", X"FEBF", X"01B6", X"FFDF", X"00C0", X"01F8", X"FE3A", X"0545", X"05AC", X"04B2", X"02ED", X"0273", X"0131", X"FE56", X"FC56", X"FA74", X"FA93", X"FA6C", X"FB10", X"FBA7", X"FD09", X"FED1", X"00D6", X"00C1", X"FF58", X"0613", X"055D", X"06CE", X"02BF", X"03F3", X"0079", X"FFFB", X"04C3", X"0142", X"FF29", X"0591", X"0778", X"03D5", X"032F", X"01D0", X"FF14", X"FDB3", X"FF33", X"FBDC", X"FB0C", X"FB92", X"FA37", X"FADC", X"FD1B", X"FFD1", X"FFF8", X"0042", X"023A", X"035C", X"02C2", X"06CA", X"07E6", X"03A4", X"0013", X"0207", X"0084", X"00ED", X"FF47", X"010C", X"01EB", X"FFD9", X"01AB", X"FF32", X"0059", X"FF55", X"0075", X"FD37", X"FD9E", X"FB7C", X"FAD0", X"FDF1", X"FF23", X"FF13", X"00D0", X"029D", X"00AE", X"005E", X"03B0", X"0437", X"0808", X"011E", X"FF74", X"FF84", X"FE52", X"0037", X"FC8F", X"FF84", X"FE6E", X"FADC", X"FCDF", X"FD2E", X"FE53", X"FE7B", X"FD6E", X"FE17", X"FB54", X"F7F0", X"FAF0", X"0017", X"FF4E", X"00D7", X"01E7", X"0075", X"00E9", X"0146", X"016B", X"04FF", X"05F6", X"01CE", X"FF6A", X"FE96", X"FEA5", X"FCF4", X"FD0D", X"FFB2", X"FBF8", X"FA50", X"FC2A", X"FC01", X"FD20", X"FBFA", X"FB2E", X"FCAC", X"FA6A", X"F8E6", X"0002", X"00B8", X"0239", X"FE69", X"FDB7", X"FE42", X"FE4B", X"FDDA", X"FFDD", X"06EC", X"066D", X"046A", X"FE97", X"FFFA", X"FD78", X"FD9D", X"FED2", X"FC84", X"F9B6", X"F7F7", X"F8E8", X"FA3E", X"FC09", X"FD39", X"FD99", X"0070", X"00A5", X"FD02", X"00F5", X"01EF", X"FE2B", X"FBC0", X"FC24", X"FA61", X"F90D", X"FBDD", X"FF57", X"039E", X"041D", X"FF3D", X"FEF7", X"004E", X"FE33", X"FD9C", X"FD31", X"F871", X"F92C", X"FAB2", X"FB5B", X"FCDC", X"FD5F", X"018C", X"0650", X"0A52", X"04B5", X"FE5D", X"FCE8", X"FEA5", X"FBAA", X"FAAD", X"FC03", X"F828", X"F75A", X"F8E6", X"F905", X"FE3F", X"FDAC", X"FDAB", X"FCA2", X"015E", X"FE53", X"FCB1", X"FDE5", X"FA67", X"FD0A", X"FDFA", X"FF96", X"003C", X"01D2", X"0546", X"0A69", X"0CC4", X"021F", X"FD7F", X"FDB7", X"FCAF", X"FD55", X"FD53", X"FC64", X"FC05", X"FB3D", X"FB05", X"FE06", X"FF94", X"FE41", X"FD9C", X"001F", X"012D", X"FE95", X"FC7C", X"020E", X"FF8B", X"017F", X"0225", X"0342", X"05A5", X"073A", X"0837", X"0A26", X"070B", X"006A", X"FD37", X"FD3A", X"FF7D", X"007B", X"FFCE", X"0058", X"FF42", X"FF23", X"FF7B", X"00D5", X"0435", X"02D4", X"FFDB", X"0091", X"01BD", X"FFCB", X"04C6", X"03EF", X"01B7", X"02C7", X"03E1", X"05BF", X"0653", X"096C", X"06A8", X"04C5", X"017B", X"FF61", X"FEBE", X"004B", X"00BC", X"018A", X"007B", X"02C5", X"02F1", X"040E", X"031B", X"04B2", X"075E", X"0706", X"0516", X"0196", X"00B2", X"01CE", X"01B2", X"05C2", X"03F3", X"02B1", X"05D5", X"04EF", X"0786", X"091D", X"044F", X"0027", X"FF36", X"FEFF", X"FFBB", X"00D1", X"0157", X"018D", X"0289", X"0402", X"0338", X"0628", X"031C", X"07A2", X"0A95", X"0A72", X"03DB", X"00D6", X"000A", X"0115", X"03C5", X"04CE", X"0565", X"05BA", X"074F", X"071E", X"0456", X"025B", X"FE90", X"FD33", X"FCCA", X"FB64", X"FDD8", X"0169", X"031E", X"0313", X"0398", X"01DE", X"0254", X"05B0", X"05EA", X"0939", X"08B3", X"0801", X"0323", X"02BF", X"FCA1", X"FFB8", X"013A", X"0563", X"0754", X"08C4", X"09D7", X"0712", X"0355", X"FE7A", X"FD03", X"FC66", X"FDCF", X"FEFD", X"FF0A", X"0089", X"0196", X"028F", X"026F", X"01E1", X"00E8", X"04CF", X"064E", X"07D7", X"0914", X"0350", X"FDEC", X"FFB4", X"FFB1", X"0159", X"FEA6", X"08A9", X"0AE4", X"0B11", X"0796", X"024E", X"000E", X"FDEE", X"FBD9", X"FE8C", X"FE2E", X"FEC5", X"010C", X"0109", X"028D", X"0206", X"0198", X"FD39", X"01AD", X"0273", X"0532", X"0218", X"020F", X"0239", X"0012", X"FF27", X"0069", X"0315", X"0402", X"0C2E", X"0D59", X"07FC", X"0492", X"01B6", X"0185", X"002C", X"FD9D", X"FFD6", X"0253", X"FE31", X"00E0", X"01EF", X"004E", X"01EC", X"021D", X"FFC5", X"FFAD", X"0263", X"0312", X"012A", X"FFB9", X"FFB9", X"0103", X"FFE6", X"FFF6", X"00DC", X"04D7", X"0973", X"0A3D", X"03F3", X"0005", X"0059", X"016F", X"006E", X"FECF", X"010A", X"015F", X"0174", X"FEB3", X"0192", X"00C6", X"004D", X"0135", X"0079", X"0154", X"00F4", X"021D", X"029E", X"FF6D", X"FEDC", X"020A", X"FF45", X"012E", X"0139", X"046C", X"06A9", X"0610", X"FF7F", X"FDD9", X"FEF9", X"FFBD", X"00E0", X"00F2", X"00FC", X"FFCF", X"0124", X"FE8F", X"0059", X"004D", X"01E8", X"01FC", X"01CF", X"012D", X"0293", X"FF6B", X"FE65", X"FFF8", X"0153", X"00F8", X"0229", X"00CA", X"0068", X"0759", X"0702", X"0560", X"0120", X"011B", X"FF82", X"FD68", X"FFFD", X"FFCC", X"FF47", X"FE00", X"FF00", X"00D3", X"FE07", X"FF02", X"FD6C", X"00C8", X"00C9", X"FEC6", X"FF63", X"FB3D", X"FBCC", X"FD29", X"0255", X"009A", X"0020", X"FFD2", X"FEBB", X"0035", X"0563", X"00EA", X"FEEB", X"FC8B", X"FC80", X"FCB9", X"FDE1", X"FCF5", X"FF6D", X"00EE", X"001D", X"0082", X"FFE8", X"FEFA", X"FF16", X"FF4A", X"FF2C", X"FD74", X"FB7D", X"FCE4", X"FAFB", X"FE45", X"010F", X"0220", X"00AF", X"FFC5", X"FE3F", X"007E", X"025D", X"013C", X"FCA5", X"F977", X"F8DF", X"F7BB", X"F99C", X"FC96", X"000A", X"FF52", X"001B", X"FFA5", X"0101", X"FFE7", X"FD25", X"FE53", X"FCDB", X"FB7D", X"FBAE", X"FD1D", X"FFD3", X"015A", X"FFD8", X"0275", X"0124", X"FEB2", X"FF3A", X"FE45", X"FE99", X"FD78", X"FAE9", X"F986", X"F58F", X"F43F", X"F441", X"F820", X"F6B5", X"F979", X"F8DE", X"F3AF", X"F8CD", X"FCAF", X"FAF8", X"FB13", X"FC5C", X"FC0E", X"FB6F", X"FC26", X"FF29", X"FEE0", X"FFA6", X"0134", X"0039", X"FFA2", X"0064", X"FF89", X"00AA", X"0024", X"FF2C", X"FCF9", X"FDC4", X"FC9B", X"FB13", X"FD4E", X"0071", X"00B9", X"FD01", X"F96F", X"FB73", X"F9C5", X"FA82", X"FAC9", X"F9FF", X"FE7A", X"FB2B", X"FAEF", X"FEDA", X"0014", X"0023", X"FF85", X"FF00"),
--        (X"00E5", X"FF48", X"018A", X"006B", X"0090", X"0034", X"FF64", X"FF45", X"00BE", X"00D5", X"FF1C", X"00A6", X"01AC", X"0168", X"013A", X"0177", X"0244", X"FFD7", X"0053", X"0153", X"00B1", X"0033", X"0054", X"FF9D", X"00BB", X"00F1", X"0128", X"00D4", X"0095", X"FF67", X"0155", X"0066", X"00D0", X"00A6", X"02B7", X"0218", X"01A6", X"039F", X"02A4", X"05BC", X"05F4", X"041E", X"0283", X"047A", X"063D", X"0574", X"0282", X"01D3", X"03D9", X"0301", X"0364", X"0232", X"00DA", X"0074", X"0175", X"0048", X"FEEF", X"00CF", X"FFFA", X"010F", X"01DB", X"021D", X"0172", X"04AA", X"0480", X"06EB", X"097A", X"0826", X"0798", X"06EC", X"06E5", X"0689", X"05D5", X"0428", X"0480", X"05D1", X"0453", X"04BF", X"03C4", X"053B", X"0109", X"0083", X"013B", X"FED1", X"FF9D", X"00AE", X"FE7F", X"0186", X"025D", X"022F", X"02E2", X"0636", X"08E9", X"0925", X"0899", X"0924", X"0ADB", X"0B61", X"09B0", X"0921", X"07F3", X"05C9", X"059A", X"05A2", X"04E9", X"03B4", X"047D", X"032D", X"06E2", X"01F9", X"00A0", X"007E", X"018A", X"FEC5", X"FE09", X"FF7C", X"FF68", X"00A0", X"0485", X"047B", X"057C", X"061B", X"05E1", X"04A3", X"0532", X"0651", X"073F", X"05CE", X"0379", X"032B", X"016F", X"FDC9", X"FDD1", X"FC84", X"FDF8", X"FFCB", X"03A0", X"06EA", X"04CE", X"032A", X"00DA", X"0057", X"FFCB", X"FF2A", X"0174", X"FD58", X"FDC9", X"00AD", X"FEAD", X"FF63", X"02ED", X"019B", X"027A", X"0436", X"0118", X"015C", X"01B3", X"04C9", X"02CD", X"02A6", X"0238", X"FF72", X"FC94", X"FB3C", X"FE47", X"0643", X"0468", X"028D", X"014A", X"016F", X"FFB7", X"FDC0", X"FFEA", X"FD61", X"FCF9", X"FDD1", X"FF8E", X"01CB", X"FF63", X"0022", X"0200", X"01F5", X"03B1", X"03C5", X"0270", X"012B", X"01FE", X"017A", X"0252", X"0095", X"FBD7", X"FD24", X"FD19", X"0423", X"01A2", X"028B", X"FEF2", X"FF11", X"FB93", X"F7FF", X"FF05", X"FF47", X"FE38", X"FD31", X"0070", X"FFE5", X"FF42", X"01A5", X"FFE2", X"021D", X"03CA", X"05B7", X"030E", X"FF3C", X"0020", X"FEAC", X"FE21", X"0132", X"FCA0", X"FE3D", X"00D4", X"04C4", X"FD86", X"0359", X"0174", X"FCD6", X"F95D", X"F7E2", X"FDA7", X"FD53", X"FF40", X"FDA3", X"FFA9", X"0075", X"017B", X"0150", X"00A6", X"00F4", X"01CA", X"015F", X"FFB9", X"FB84", X"FCC1", X"FEEC", X"00D5", X"FFAA", X"FDEA", X"002C", X"04CA", X"0429", X"035C", X"034C", X"FF3B", X"FCBE", X"FB7C", X"FB49", X"FE2E", X"FF70", X"FEB6", X"FFC6", X"014D", X"00F1", X"02DE", X"0123", X"019B", X"013A", X"014D", X"FE35", X"FE3F", X"FCE4", X"FEAC", X"FEDA", X"001B", X"0057", X"FF6D", X"0255", X"03A1", X"051F", X"0638", X"FFD9", X"FEBC", X"FB34", X"FCC0", X"FF73", X"FE21", X"FF49", X"0199", X"02EE", X"00AE", X"00D7", X"011C", X"016C", X"014E", X"0335", X"FFEF", X"F9D0", X"FB6B", X"FD11", X"FEDC", X"FF16", X"FEDB", X"FE4D", X"002D", X"03F7", X"0954", X"06DC", X"068B", X"0017", X"FFD1", X"FC33", X"FC1B", X"FD7C", X"FDAF", X"0207", X"0265", X"0119", X"FF24", X"FEC2", X"FEC8", X"FF5A", X"01EC", X"02EB", X"FCE6", X"F8BA", X"FAE3", X"FB42", X"FD55", X"FF13", X"FF44", X"FDE1", X"0199", X"0715", X"0AE9", X"082C", X"03AA", X"FEE4", X"006D", X"FC96", X"FB1E", X"FDFA", X"FE7C", X"022A", X"0086", X"FD8D", X"FC63", X"FE0C", X"FDF8", X"FE0F", X"02A6", X"034B", X"FB45", X"F9FE", X"F91C", X"FDD3", X"FC39", X"FDBB", X"0054", X"00D0", X"01CB", X"0536", X"061A", X"031F", X"0250", X"FDEA", X"FF8D", X"FF3B", X"FA7A", X"FD15", X"FCD6", X"001F", X"FE5D", X"FB6C", X"FD4C", X"FDA8", X"FF24", X"0264", X"041C", X"00BA", X"FB26", X"FB49", X"FCC3", X"FDFD", X"FD3D", X"FD04", X"FE03", X"FDE6", X"00DB", X"0602", X"0476", X"03A6", X"03E9", X"0241", X"0098", X"FDB9", X"FA96", X"FB88", X"FB4B", X"FC51", X"FD91", X"FCE6", X"FBCE", X"0090", X"035F", X"025C", X"03D6", X"FFE9", X"FC1B", X"FC39", X"FE2C", X"FBFD", X"FB4C", X"FC16", X"FE1D", X"0022", X"005F", X"0141", X"03A2", X"037F", X"0630", X"01DD", X"FFD6", X"FFC1", X"FB91", X"FC37", X"FC79", X"FF88", X"FFF1", X"FDC5", X"FDB0", X"006C", X"0325", X"0363", X"0236", X"FE7D", X"FC48", X"FD81", X"FD80", X"FBB9", X"FBC3", X"FCB2", X"FDAA", X"FF36", X"0013", X"0179", X"07FF", X"0682", X"0464", X"02A0", X"FEC7", X"FFAF", X"0158", X"FFF7", X"FE98", X"023F", X"001D", X"FD40", X"FD2F", X"00B9", X"02F3", X"02BD", X"0111", X"FD7B", X"FC89", X"FB7B", X"FDE2", X"FC35", X"FE46", X"FF76", X"FF16", X"FDA4", X"032A", X"0451", X"0854", X"0A13", X"0996", X"03A6", X"FFC2", X"FEFA", X"FF99", X"02B4", X"010D", X"0369", X"05F9", X"0468", X"04AB", X"038B", X"05C4", X"04A3", X"0229", X"FFAF", X"FD80", X"FE2B", X"009E", X"00AA", X"02A6", X"022B", X"0234", X"019A", X"0554", X"061B", X"09AD", X"08D7", X"0452", X"023C", X"0037", X"FDCB", X"0027", X"015B", X"04AF", X"0740", X"0A90", X"08B4", X"0619", X"0747", X"08F2", X"073F", X"0279", X"FF1B", X"FFA6", X"01CD", X"03AB", X"0642", X"06A4", X"077B", X"03B8", X"05DA", X"096A", X"0AE2", X"0B5D", X"07B2", X"FEC4", X"FE63", X"FEA4", X"FEBB", X"0079", X"018A", X"0540", X"0A71", X"09B0", X"0793", X"07A1", X"0754", X"07E2", X"06CA", X"0563", X"030F", X"0043", X"0224", X"0640", X"05EB", X"0876", X"07CC", X"0663", X"0628", X"0CAB", X"0CBD", X"0972", X"0575", X"0296", X"FD2F", X"FFCD", X"0183", X"04A5", X"0853", X"086A", X"0500", X"058A", X"0646", X"05EC", X"05C7", X"0538", X"03E9", X"042B", X"029F", X"FF70", X"02EC", X"0258", X"0571", X"0717", X"0766", X"08BD", X"0769", X"08E0", X"093E", X"0A3B", X"0536", X"0206", X"FF48", X"0132", X"01A9", X"04D2", X"07C9", X"02A0", X"FF36", X"FFDE", X"01A8", X"0101", X"0237", X"FEDA", X"01FD", X"02B7", X"0543", X"0327", X"011D", X"00FB", X"0320", X"0413", X"03EE", X"0509", X"04BF", X"06BF", X"05E5", X"045A", X"02D2", X"02B8", X"FFC7", X"002C", X"FEB8", X"02C6", X"05E5", X"0005", X"FA57", X"FC7A", X"FBBF", X"FDD6", X"FD8D", X"FC73", X"01BF", X"02DF", X"0327", X"0271", X"FF71", X"0063", X"FF37", X"01D8", X"02C4", X"0527", X"042C", X"04AE", X"04D8", X"027F", X"FEE4", X"FE33", X"0026", X"FFEC", X"FF99", X"03D4", X"0840", X"FC62", X"F9DB", X"F832", X"FADA", X"FCE5", X"FD01", X"FDB9", X"00EF", X"020A", X"0158", X"00E7", X"FF99", X"FFB0", X"FFE0", X"01FF", X"03C7", X"03DE", X"0630", X"0255", X"05D4", X"01B4", X"FDDD", X"FC63", X"010D", X"FF0B", X"FF58", X"00ED", X"0294", X"FDBC", X"F7BE", X"FB1A", X"FC4B", X"FE7E", X"0048", X"007E", X"01FC", X"0297", X"0249", X"034F", X"0335", X"05A8", X"03B3", X"0246", X"01C3", X"0255", X"024B", X"037E", X"044A", X"04F8", X"00BC", X"0050", X"FE8E", X"FF6E", X"0049", X"034B", X"FE5D", X"FB58", X"FBE8", X"FE3D", X"FC6A", X"FD56", X"00D1", X"FFCE", X"0142", X"00F3", X"0194", X"016D", X"0293", X"0346", X"0396", X"03CA", X"02CD", X"032C", X"0348", X"0094", X"FF3F", X"FFFA", X"FE5E", X"003B", X"0088", X"FFE9", X"FF00", X"005E", X"00AD", X"0142", X"004E", X"FE53", X"FCFF", X"FCAC", X"FE1F", X"FD7D", X"020E", X"FFA4", X"00D8", X"FD4D", X"FC4D", X"FBF0", X"FE03", X"FEC5", X"FC6E", X"025B", X"0170", X"00C4", X"0164", X"0015", X"001C", X"FF1B", X"FEB2", X"00F9", X"FFA5", X"0059", X"0044", X"FE31", X"FF82", X"FFAE", X"FF16", X"FDA2", X"FC80", X"FDF6", X"00CD", X"FF0D", X"FBA6", X"F9E3", X"FA3C", X"FCEF", X"FB88", X"FB8B", X"FB9E", X"FEEE", X"FC72", X"FDC1", X"FEA0", X"000A", X"00D6", X"00DF", X"FFEF"),
--        (X"015C", X"0123", X"0225", X"00DC", X"FE8E", X"FFAA", X"015B", X"FF95", X"005F", X"005C", X"0008", X"FF8A", X"0142", X"006F", X"0042", X"004B", X"009F", X"0069", X"FF85", X"FF37", X"0095", X"002B", X"0061", X"0265", X"FFC7", X"FF53", X"FEBE", X"FE64", X"FE66", X"FF57", X"01E8", X"0124", X"FF14", X"FFD5", X"00B0", X"0274", X"03A6", X"02D7", X"032D", X"0542", X"0493", X"03D9", X"0129", X"0514", X"0493", X"0537", X"0333", X"039C", X"030F", X"046C", X"026A", X"030D", X"018F", X"FFDB", X"0063", X"0142", X"0058", X"017E", X"00D9", X"0152", X"00E9", X"0018", X"040F", X"05C6", X"0657", X"0793", X"0A9A", X"0C4C", X"0983", X"0AE8", X"0B33", X"0A5D", X"09AC", X"06D9", X"05CB", X"07E6", X"0589", X"06A5", X"0400", X"03E3", X"0376", X"02E9", X"01E8", X"018D", X"00FA", X"0165", X"FD67", X"024F", X"03FB", X"0113", X"04DF", X"078C", X"0B13", X"0AEE", X"0A1B", X"0A14", X"09DB", X"08A4", X"0723", X"050C", X"019E", X"0323", X"FFBF", X"045F", X"06E4", X"0445", X"026C", X"FF15", X"FF89", X"0172", X"0164", X"FF10", X"012E", X"003F", X"FDAB", X"FF92", X"FCDB", X"FEFD", X"FF80", X"FF88", X"FE45", X"018E", X"FE50", X"FE5E", X"FE36", X"FE94", X"FDC5", X"0015", X"0020", X"014A", X"FDCF", X"FDDD", X"FE32", X"0066", X"00AB", X"0449", X"03D8", X"0132", X"014C", X"00F2", X"FFA8", X"0079", X"FE50", X"FE02", X"FCFC", X"F9E3", X"FC8B", X"FF16", X"004C", X"0070", X"FF96", X"FE9F", X"FCBB", X"FE25", X"FFE5", X"FE0A", X"FFCF", X"0099", X"00E5", X"00DC", X"FFD8", X"FF17", X"0037", X"00F8", X"008C", X"00F0", X"0155", X"018E", X"FE9E", X"FE96", X"022C", X"FCE4", X"FBA9", X"FCE2", X"FDFE", X"FF96", X"FD3F", X"FDEA", X"FF47", X"0017", X"FEA9", X"001E", X"01A5", X"0214", X"000F", X"FFEF", X"0067", X"022B", X"FFE1", X"FF61", X"00B6", X"FF3E", X"01EE", X"FED4", X"FF51", X"0179", X"007A", X"FBEF", X"0087", X"FA1A", X"F871", X"FE42", X"FEE1", X"FE64", X"FDAB", X"FEC8", X"00A2", X"02B5", X"0177", X"022A", X"0309", X"00D3", X"FF34", X"00E5", X"00C3", X"0041", X"000F", X"0018", X"FF6B", X"010E", X"022A", X"0246", X"FE28", X"01CA", X"0333", X"FFE3", X"0046", X"F8AF", X"F6D2", X"FD0A", X"FDA5", X"FECB", X"0004", X"FFC1", X"00B5", X"0257", X"0055", X"00A4", X"0317", X"0150", X"FF88", X"FEFC", X"FD66", X"FE87", X"FFB2", X"0025", X"FF28", X"0631", X"05AD", X"0346", X"FF72", X"FF35", X"FF8C", X"FE22", X"FE7F", X"F894", X"FA24", X"FD44", X"FDF7", X"FEC5", X"0085", X"014A", X"013E", X"018F", X"0131", X"00FA", X"FEF7", X"FC6A", X"FAE2", X"FD07", X"FAAD", X"FCD9", X"FDAC", X"FE31", X"00E6", X"069B", X"0BE3", X"07AC", X"0223", X"01FB", X"FFAC", X"FE55", X"FE04", X"FBCA", X"FF3D", X"00BA", X"00E4", X"0206", X"022B", X"0399", X"015D", X"035E", X"016A", X"019D", X"021F", X"FBCF", X"FB5A", X"FBD6", X"FD13", X"FBA1", X"FB4C", X"FBA8", X"FDFC", X"07A0", X"0E4E", X"0B6F", X"0632", X"FDFF", X"0042", X"0047", X"FBB7", X"FB78", X"0079", X"00E3", X"0031", X"0180", X"024C", X"0070", X"FE05", X"FF32", X"FE59", X"01BC", X"FBCB", X"F928", X"FC9C", X"FC95", X"FBA1", X"FBAF", X"F986", X"FB39", X"FA4B", X"024E", X"085D", X"08BB", X"0120", X"FFD4", X"FFC1", X"FEF3", X"FB17", X"FE10", X"FEA8", X"FE5E", X"FF9D", X"FE69", X"FEF1", X"FF17", X"FFA1", X"0055", X"00AB", X"FE8A", X"FAD3", X"F81C", X"F870", X"FA03", X"FC0A", X"F951", X"F8BF", X"F874", X"F88B", X"F9F5", X"0052", X"01E2", X"0213", X"0268", X"014B", X"FF4A", X"FE9B", X"FEDE", X"FDE3", X"FE46", X"005F", X"FF53", X"FE25", X"FF1B", X"FFBF", X"011A", X"007C", X"FD74", X"FACF", X"F834", X"F838", X"FACC", X"FA4B", X"FAB7", X"FA98", X"FC52", X"FCE5", X"FE7B", X"0305", X"FEE6", X"05C1", X"0148", X"036D", X"FEDF", X"FD88", X"FC36", X"FCC9", X"00A7", X"014D", X"00D3", X"FE9D", X"017D", X"024B", X"006E", X"FEA4", X"FB96", X"FAFC", X"F8DE", X"F7B5", X"F9B5", X"FA5F", X"FCEE", X"0073", X"010D", X"0158", X"03DD", X"05F9", X"02DA", X"03F9", X"0176", X"00DA", X"FF5B", X"FDB8", X"FC38", X"FCC4", X"0110", X"0315", X"0112", X"018D", X"0221", X"0300", X"0172", X"FE57", X"FA41", X"F88C", X"F8B6", X"FB13", X"FBF5", X"FE90", X"0179", X"01F1", X"0209", X"022E", X"0393", X"079E", X"04AE", X"0194", X"01A4", X"FCC2", X"FC79", X"FD51", X"FC3D", X"FD0F", X"01C9", X"02AF", X"FEA9", X"FBFF", X"FE43", X"00DA", X"01DF", X"FE38", X"FABF", X"F9E9", X"FABC", X"FCBC", X"0108", X"0437", X"0523", X"02CB", X"037A", X"0453", X"03E6", X"05C8", X"0822", X"047F", X"0333", X"00A0", X"FDBD", X"FEBF", X"FC61", X"FF02", X"05E4", X"06C5", X"0072", X"FD4D", X"FED0", X"0389", X"0051", X"FD0A", X"FB13", X"FC66", X"010E", X"01B7", X"04AC", X"0527", X"048A", X"04C4", X"037C", X"0362", X"0437", X"05EE", X"0A47", X"03A5", X"03B7", X"FE04", X"FF30", X"FC9F", X"FA24", X"FF31", X"0421", X"058F", X"0328", X"00E8", X"006E", X"0459", X"03BA", X"0397", X"020C", X"021B", X"0351", X"05A1", X"0529", X"0520", X"047B", X"023C", X"0346", X"04B3", X"088D", X"0B5A", X"09C6", X"FEAB", X"00E9", X"FFF6", X"009F", X"FFE3", X"FC3D", X"00E1", X"01E4", X"02B5", X"0407", X"0536", X"04FF", X"0351", X"096E", X"088D", X"06C4", X"04A3", X"052A", X"02D9", X"0364", X"0494", X"049C", X"0395", X"02E1", X"0553", X"05CC", X"0947", X"07D3", X"00EC", X"FF23", X"FE41", X"01B6", X"FDF4", X"FF27", X"007B", X"0320", X"FFE0", X"0026", X"034F", X"03EC", X"0612", X"069E", X"03F6", X"02A4", X"01DB", X"00E7", X"02D1", X"03A1", X"0369", X"037C", X"029D", X"036C", X"04FB", X"0565", X"06DC", X"0799", X"00D0", X"004E", X"0108", X"0072", X"FF83", X"01B8", X"019E", X"0029", X"FF10", X"0110", X"0128", X"04A4", X"0238", X"020F", X"0191", X"0027", X"0045", X"0089", X"FF44", X"00E5", X"00EF", X"0202", X"02D9", X"0563", X"05CB", X"0976", X"066C", X"05A5", X"0435", X"006C", X"FEF0", X"FF9D", X"FDC8", X"00FD", X"000A", X"FFCC", X"FFE1", X"0034", X"01B6", X"00D0", X"0111", X"001A", X"0149", X"FFBE", X"FF88", X"FDDD", X"FEE9", X"FD7E", X"FF3C", X"008A", X"0078", X"02AF", X"0398", X"0543", X"0407", X"0586", X"0286", X"007E", X"00FB", X"FFFA", X"FEDD", X"FFA9", X"00DD", X"01A5", X"0185", X"FFFE", X"0254", X"024D", X"02D9", X"00B4", X"010D", X"FD7D", X"FDB0", X"FD97", X"FE4A", X"FD05", X"FA45", X"FCDB", X"FE6B", X"FEFD", X"0093", X"0004", X"FF7A", X"0150", X"011F", X"0039", X"FFCD", X"FEED", X"FCE4", X"0090", X"FD0F", X"FE18", X"00A6", X"0179", X"0253", X"0464", X"013A", X"0130", X"0332", X"0306", X"02F4", X"0111", X"00C8", X"01FB", X"FFAC", X"FE73", X"FD69", X"FEE0", X"FE51", X"FC96", X"03B6", X"03C6", X"0387", X"FD95", X"FF6C", X"FF1F", X"FF5B", X"016F", X"FF7B", X"FCCD", X"FE47", X"FE3C", X"FEDB", X"FFC9", X"FF8C", X"0090", X"00EA", X"0248", X"FFF3", X"0296", X"02AE", X"02BE", X"0174", X"002A", X"FCD4", X"FE04", X"0136", X"020E", X"018A", X"0273", X"01CF", X"FF10", X"FFDA", X"0093", X"FF8E", X"00FB", X"FF09", X"FD47", X"FC28", X"F7B8", X"F6FB", X"FB98", X"FD82", X"FFF3", X"019B", X"00B7", X"FE30", X"03D8", X"FF8F", X"FE8A", X"FDFF", X"0009", X"FE72", X"FE7C", X"FF89", X"FC76", X"FD2C", X"FFCC", X"0093", X"FF81", X"0100", X"FF88", X"FF95", X"0087", X"0027", X"00F8", X"006E", X"001C", X"FF08", X"FE96", X"01A0", X"0286", X"011E", X"003F", X"FB01", X"FCC8", X"FD43", X"FD35", X"FC8A", X"FC72", X"FDC4", X"FA35", X"FAF5", X"FCD7", X"00FD", X"0070", X"005F", X"00E5"),
--        (X"FED2", X"0026", X"FF42", X"FFB0", X"00D8", X"FF56", X"FFF8", X"FF15", X"00BB", X"00EC", X"004E", X"FFFD", X"FFF0", X"FFC7", X"00C0", X"00A1", X"0164", X"0098", X"0076", X"FFB9", X"0088", X"01A9", X"FF1B", X"FED1", X"FF01", X"00D1", X"FE83", X"FFE0", X"0107", X"FEA3", X"FFFC", X"FF07", X"001B", X"0014", X"006E", X"FD9C", X"FF64", X"FC54", X"FEC7", X"0077", X"FD3C", X"FDF5", X"015D", X"0296", X"02B1", X"0241", X"FE79", X"FF6C", X"FDC2", X"FF29", X"00CC", X"FFD3", X"00C9", X"0001", X"0032", X"FFBD", X"FF39", X"FFAA", X"006B", X"00E3", X"FF25", X"FE9A", X"FCA8", X"FD84", X"FD0C", X"FE1D", X"FE2E", X"FA8B", X"FDCE", X"001C", X"01C5", X"0123", X"0319", X"012B", X"FF9E", X"FE84", X"FE42", X"FD5A", X"FC16", X"FE51", X"00B8", X"0236", X"FF10", X"FFCD", X"00AE", X"FF7C", X"02DD", X"027C", X"FE56", X"FCF7", X"FC81", X"FDD0", X"0100", X"011E", X"FF8B", X"001D", X"0286", X"03DC", X"014F", X"0096", X"0079", X"0161", X"FD92", X"FDE1", X"FEB1", X"FB02", X"F9A4", X"FC29", X"FD07", X"00E8", X"FE34", X"012D", X"FF4D", X"0072", X"0252", X"015B", X"FDBD", X"FD35", X"014F", X"02CA", X"04E4", X"044E", X"0476", X"07F1", X"05EA", X"0866", X"05A1", X"05A0", X"03AE", X"0350", X"01AA", X"FE61", X"FC3D", X"FBDC", X"FB3D", X"F9CF", X"FA01", X"FEC4", X"0256", X"FF5A", X"003A", X"FFF4", X"026D", X"0127", X"FEFB", X"001B", X"01C9", X"0119", X"FE68", X"0071", X"0312", X"04E0", X"01E0", X"02F0", X"02ED", X"02F6", X"0481", X"0390", X"00FD", X"00D9", X"FDF5", X"FE20", X"FCDE", X"F897", X"FA2B", X"FF60", X"FE95", X"FDCE", X"FF33", X"00F7", X"FF23", X"FF4F", X"FF14", X"FD5B", X"FE8C", X"FC0C", X"FE6D", X"FD3F", X"0117", X"01E8", X"0162", X"0181", X"FFE2", X"00E1", X"0192", X"FF78", X"00FA", X"025B", X"0114", X"00D4", X"0035", X"FCF2", X"FCF9", X"FC73", X"FCEC", X"FC8C", X"00F0", X"FED9", X"FC86", X"FD0D", X"FE47", X"FDD3", X"FF14", X"FF15", X"FE1B", X"FE03", X"FFF3", X"00D5", X"0128", X"0269", X"01D9", X"0085", X"0201", X"010F", X"03D9", X"0232", X"0250", X"01D4", X"0387", X"0297", X"FDD3", X"FDF3", X"FDEC", X"FE7A", X"0192", X"FE10", X"FC58", X"FE48", X"FF7A", X"0076", X"0068", X"FE10", X"FED5", X"FFB1", X"00D8", X"FF1E", X"02F1", X"033A", X"00DA", X"0153", X"0257", X"0152", X"03E8", X"04D6", X"0425", X"04F3", X"0507", X"04A5", X"03D8", X"FE6E", X"02A6", X"043A", X"0060", X"FB90", X"FE37", X"0049", X"0105", X"004D", X"FFF4", X"0084", X"0085", X"FE3E", X"0155", X"005F", X"0189", X"00DF", X"0168", X"025F", X"0388", X"05BC", X"03E1", X"047A", X"0485", X"0405", X"055B", X"06F6", X"06FA", X"04A0", X"00CE", X"FD9A", X"FD60", X"FA12", X"FE1A", X"FEE2", X"0148", X"FFB8", X"FF97", X"FF84", X"FE8F", X"FE4D", X"FF42", X"FFC5", X"0069", X"FFA4", X"02AF", X"0114", X"021B", X"0251", X"032A", X"02C3", X"0423", X"0507", X"0356", X"06FC", X"0835", X"03DA", X"022A", X"FFB7", X"FEE1", X"FFAD", X"FE6E", X"FDA6", X"007E", X"00B0", X"FEA1", X"FE5D", X"FD5B", X"FD55", X"FD88", X"FDAC", X"FB85", X"FF39", X"0151", X"FE63", X"FCD4", X"FDE2", X"FF94", X"0258", X"00D5", X"FF0F", X"008C", X"0701", X"08EF", X"0769", X"0657", X"026C", X"FE9A", X"FD49", X"FAF7", X"FE0D", X"FEC6", X"FEF1", X"FE0C", X"FE9B", X"FD5A", X"FC90", X"FC6A", X"FA9A", X"FD23", X"FF5A", X"014C", X"FD8C", X"FBC7", X"FACF", X"FE5B", X"00D5", X"0192", X"0013", X"FF5E", X"0011", X"0745", X"04EF", X"0621", X"02A4", X"01B1", X"FFB8", X"FC98", X"0134", X"FCEB", X"FC03", X"FCE8", X"FEA2", X"FF3C", X"FF38", X"FC57", X"FC45", X"FDA7", X"0224", X"006A", X"FD9C", X"FB12", X"FC34", X"FE83", X"FFF7", X"FF95", X"FB8E", X"FA4B", X"FE8A", X"FFA8", X"02F8", X"03DC", X"02A2", X"0016", X"FDA4", X"FD50", X"FF35", X"FE54", X"FAD3", X"FDD6", X"FEE0", X"FFB7", X"FF46", X"FD1F", X"FB6A", X"FFD4", X"0256", X"02FC", X"FE94", X"FBEA", X"FB4A", X"FE43", X"FB21", X"FAEA", X"FAE7", X"FA0D", X"FC55", X"FF0D", X"FE1A", X"0538", X"0188", X"003F", X"FEBC", X"0284", X"0129", X"02BE", X"FF68", X"FCDE", X"FE8E", X"FEF9", X"0046", X"FE3F", X"FCDA", X"004F", X"04E9", X"032E", X"FC8E", X"FB00", X"FA2A", X"FA23", X"FB0C", X"FA2E", X"FAF2", X"F902", X"FE05", X"01A0", X"00E7", X"04CC", X"03D9", X"FEAA", X"FFBD", X"0426", X"05A3", X"052B", X"0415", X"FE92", X"FCFA", X"FD57", X"FEBE", X"FDBC", X"FBCA", X"03C3", X"043A", X"FFCC", X"FC96", X"FB6C", X"FAAD", X"F929", X"FB0F", X"FCC4", X"FE0D", X"0060", X"01C2", X"0263", X"02B0", X"0441", X"02ED", X"0060", X"020D", X"0265", X"05DB", X"06C3", X"0658", X"024F", X"FC44", X"FA22", X"FC89", X"FBC3", X"FDE8", X"0100", X"FF9F", X"FF56", X"FBE7", X"FCB2", X"FB50", X"FAD7", X"FDF5", X"0116", X"0068", X"02C2", X"04D8", X"05AC", X"015A", X"031C", X"02F8", X"FDDF", X"0051", X"01B3", X"03B5", X"05C0", X"0639", X"050F", X"01EC", X"000D", X"FBD9", X"FE06", X"FC90", X"FE0A", X"FED8", X"FDD9", X"FD5C", X"FE60", X"FE72", X"FEDA", X"00C5", X"028B", X"0234", X"0866", X"07C1", X"0690", X"04D1", X"003B", X"02A5", X"FF3A", X"0265", X"012D", X"0198", X"02BC", X"06A4", X"0581", X"03D4", X"042A", X"03BA", X"00F0", X"FC76", X"FDD8", X"FFF6", X"FE55", X"004B", X"FF41", X"0137", X"014B", X"021E", X"0411", X"0663", X"08C8", X"090B", X"0490", X"05B4", X"0439", X"0231", X"0035", X"026F", X"0217", X"035B", X"03FA", X"0707", X"0905", X"0780", X"06B6", X"0500", X"02FA", X"0120", X"FD6A", X"FEE1", X"FEEE", X"0224", X"0027", X"018D", X"0364", X"04E4", X"069E", X"0728", X"09F3", X"04F5", X"01F4", X"0252", X"029C", X"FEFA", X"000B", X"0075", X"02C7", X"03F3", X"02B6", X"0665", X"07CD", X"081C", X"02FA", X"0326", X"026C", X"01F4", X"FE93", X"FF56", X"01E6", X"012F", X"00D5", X"0321", X"0672", X"068C", X"073A", X"0814", X"0727", X"04CC", X"FFCF", X"018D", X"00D8", X"0060", X"FFE9", X"FED2", X"0493", X"036B", X"040D", X"063F", X"07F9", X"0459", X"0244", X"02CA", X"00A6", X"01A3", X"01F4", X"0273", X"0225", X"03A8", X"032A", X"04CD", X"077F", X"061C", X"06A6", X"04D8", X"052A", X"01E2", X"FE9E", X"0199", X"FFCC", X"FEFA", X"FF8B", X"0101", X"0402", X"0251", X"052C", X"0511", X"02CB", X"0262", X"01AC", X"01EE", X"007E", X"02C7", X"0395", X"03BB", X"03F2", X"041A", X"0525", X"060A", X"066C", X"038C", X"03E4", X"00F4", X"000D", X"02FF", X"FF37", X"FFBE", X"FF4C", X"FFEE", X"FFA7", X"0043", X"0122", X"0228", X"0111", X"FD52", X"FC00", X"FD1B", X"FC67", X"FE4D", X"0030", X"FE97", X"0285", X"023B", X"02B9", X"030E", X"0253", X"FFEF", X"038E", X"01F3", X"FE83", X"FDA5", X"FF25", X"FDAA", X"0472", X"02F1", X"0220", X"FF32", X"FFCC", X"0107", X"00DF", X"FFDE", X"002A", X"FCDC", X"FB58", X"FAA1", X"FD61", X"FD13", X"FDCF", X"FD87", X"FF01", X"FFAD", X"FF6E", X"FF2E", X"FFCB", X"01B8", X"003E", X"0027", X"FDB6", X"FD7C", X"FE27", X"FDC2", X"014C", X"FF8C", X"01A1", X"FFD1", X"FF9E", X"FF80", X"009D", X"FE2C", X"FCC4", X"FBDB", X"F832", X"F9D9", X"FAA2", X"F9D8", X"FCC2", X"FE0F", X"FE7D", X"FDE1", X"FD02", X"FC3B", X"FD7D", X"0011", X"FDDF", X"FFAC", X"FDC0", X"FC36", X"FC93", X"FD41", X"FEB2", X"00FD", X"FFE6", X"FFB4", X"FF9E", X"FF86", X"FF48", X"000E", X"FF92", X"FEA7", X"FEF5", X"FDF7", X"FE2F", X"FDC8", X"FC54", X"FF1F", X"FF85", X"FCBF", X"FA0C", X"FA21", X"FA7A", X"F9FE", X"FBD5", X"FA5B", X"FE06", X"FAB0", X"FC56", X"FC66", X"FFEF", X"FFA5", X"0040", X"FF87"),
--        (X"0020", X"0092", X"0033", X"FEEF", X"00A8", X"006D", X"005E", X"FE82", X"0130", X"FE51", X"FFC5", X"012D", X"0192", X"012E", X"FF2E", X"00B5", X"0164", X"0018", X"FF26", X"FF68", X"FF6F", X"FF93", X"FFE6", X"01BC", X"00A6", X"FF09", X"00FE", X"FF68", X"FED6", X"0009", X"FFD6", X"FFEA", X"001F", X"FFCF", X"0474", X"03C9", X"0384", X"031C", X"029D", X"02D6", X"0498", X"04C5", X"FE31", X"00F1", X"FEC3", X"039E", X"05E8", X"0767", X"0638", X"02EF", X"02FC", X"0097", X"FE7A", X"0065", X"00BD", X"000E", X"FEF2", X"FFA9", X"FFF5", X"0156", X"044A", X"0155", X"05BB", X"055A", X"04A3", X"FC5E", X"FC70", X"FDF9", X"FF2B", X"00D1", X"0026", X"0007", X"00BE", X"0373", X"05BF", X"079D", X"06E3", X"07CC", X"06AE", X"0535", X"02AE", X"0103", X"FF9F", X"0131", X"FEA5", X"00E5", X"003C", X"01A7", X"021A", X"01F2", X"007A", X"00C4", X"015B", X"FE7F", X"00BE", X"FEF9", X"013B", X"0180", X"0189", X"05E1", X"044A", X"05CE", X"084C", X"06AD", X"05CD", X"03BC", X"0527", X"05FD", X"06AB", X"024E", X"01A6", X"FFCC", X"FF55", X"007A", X"FE9C", X"0313", X"0212", X"FE6F", X"FBFD", X"00A3", X"FE61", X"FE58", X"FDF8", X"FE5E", X"FEA3", X"FE88", X"FE41", X"014B", X"02FA", X"0304", X"02AE", X"01B9", X"0158", X"02C6", X"0181", X"0213", X"04B4", X"0416", X"0487", X"011F", X"FF80", X"0066", X"FE6D", X"FF83", X"FDA5", X"FC73", X"FF78", X"FDCF", X"FDEA", X"FD1E", X"FE0A", X"FC70", X"FDF0", X"FEAC", X"FF3C", X"FEEA", X"01BF", X"0051", X"00FF", X"0232", X"02AC", X"032A", X"00B1", X"FFA7", X"009C", X"015F", X"047E", X"0193", X"005B", X"0147", X"FDD0", X"FE88", X"FE44", X"006D", X"FEAC", X"FD4F", X"FC2F", X"FDA2", X"FD4E", X"FE8B", X"FF7D", X"FF9A", X"016C", X"01FF", X"021A", X"01B7", X"0023", X"00C0", X"01FA", X"01DD", X"02E7", X"0291", X"02DD", X"03B7", X"00C8", X"0156", X"FF84", X"026E", X"FC40", X"FCF5", X"FF59", X"FF9D", X"FD7A", X"FD7A", X"FFF5", X"FF85", X"00EE", X"FEA5", X"0095", X"FEE0", X"01EF", X"03B5", X"02BF", X"0295", X"01FC", X"00BC", X"007C", X"0146", X"008B", X"02BD", X"03EE", X"03DD", X"FF97", X"017B", X"0190", X"FE24", X"FB15", X"FDD2", X"FFB1", X"FF1B", X"FE3F", X"FED3", X"FF9D", X"00C7", X"00C5", X"FE82", X"FDB6", X"FFF6", X"0105", X"021A", X"0423", X"02F1", X"013D", X"027E", X"0217", X"03D8", X"0210", X"0387", X"0456", X"0120", X"02D7", X"0413", X"FF85", X"FD08", X"FD92", X"FD14", X"FF60", X"FD53", X"FEA5", X"00D3", X"0203", X"00B9", X"FF25", X"FECF", X"FDBF", X"00BE", X"00E9", X"FDE4", X"0167", X"FFC8", X"FF31", X"000D", X"01E5", X"0434", X"05D3", X"04B9", X"0611", X"067A", X"07F4", X"01AA", X"FEC4", X"FCF5", X"FCE0", X"025D", X"013E", X"FFA9", X"FEB1", X"02B3", X"0293", X"019B", X"FFD3", X"FDE4", X"FF5E", X"02C0", X"043C", X"FFA4", X"FE27", X"FD23", X"FDA6", X"FF29", X"FF3D", X"0045", X"04F2", X"0A65", X"0B06", X"0756", X"05E2", X"019A", X"FEA6", X"FB0E", X"FC39", X"FE72", X"FF43", X"FEA3", X"030F", X"0214", X"0105", X"0171", X"FDB1", X"FED1", X"000A", X"0735", X"07C0", X"FDE5", X"FDAA", X"FE5A", X"FE1C", X"FB17", X"FB83", X"FE56", X"0303", X"0B8F", X"0E6A", X"0782", X"0563", X"0082", X"FF6B", X"FB86", X"F8B3", X"FE63", X"FFD7", X"03CB", X"04ED", X"043F", X"004C", X"0080", X"00E4", X"0017", X"01B8", X"079E", X"0520", X"FCFA", X"FDAF", X"00BB", X"FCE2", X"FBE4", X"FA0A", X"FC60", X"0438", X"0B7A", X"0953", X"021B", X"FE34", X"FD77", X"FEE2", X"FFD9", X"FA24", X"0020", X"FF1E", X"0289", X"0389", X"0152", X"FFE1", X"0228", X"0034", X"0177", X"05C4", X"05DC", X"0079", X"FD14", X"FCBD", X"FCDF", X"FCCA", X"F9D3", X"F859", X"FCC2", X"04A3", X"084F", X"028F", X"F8DC", X"F811", X"FC22", X"00BB", X"00CD", X"FC0D", X"FC4C", X"FA8C", X"FF26", X"0015", X"FE16", X"FC75", X"01FA", X"014E", X"054C", X"06A3", X"03C0", X"FE1A", X"FBA5", X"FC4F", X"FC6E", X"FA7F", X"F792", X"FB2A", X"0331", X"06BB", X"0090", X"FE6D", X"F7FC", X"F796", X"FC2C", X"FF0A", X"0001", X"0058", X"F9FD", X"F9A7", X"FEF4", X"FD1A", X"FDD8", X"FDCB", X"00F8", X"035C", X"06A1", X"05D1", X"FFD6", X"FB90", X"F8D6", X"FA5C", X"FAAE", X"FBA8", X"FAEF", X"FEB9", X"046C", X"0483", X"011B", X"FEA9", X"F684", X"F6A2", X"FC4C", X"FF71", X"0288", X"02FC", X"FD1F", X"FDAE", X"FDF8", X"FF03", X"FBED", X"FD5C", X"00AE", X"02CB", X"044E", X"01E0", X"FC2E", X"F96B", X"FA22", X"FA85", X"F99A", X"FD3E", X"FE16", X"0145", X"0150", X"02FC", X"014E", X"FDAA", X"F3E2", X"F52E", X"FD15", X"0086", X"02B3", X"008F", X"FE45", X"FEE0", X"FE4F", X"0223", X"FE7B", X"FFCC", X"01B7", X"018A", X"02D9", X"FE4A", X"FA02", X"F5DC", X"F8B9", X"FD4D", X"FD61", X"FF73", X"0207", X"00DE", X"00BA", X"FFBB", X"FF55", X"FBA3", X"F1F6", X"F7CF", X"0091", X"FD21", X"00D3", X"010E", X"FF20", X"FE6C", X"00C8", X"026C", X"007C", X"0083", X"0377", X"035A", X"FFE9", X"FBD7", X"FC0E", X"F898", X"FC71", X"FDDD", X"FEB0", X"012E", X"0392", X"023F", X"0047", X"0109", X"FDE3", X"FA70", X"F4A9", X"F916", X"FC0C", X"FEE8", X"0091", X"01B7", X"FF2F", X"FE16", X"0214", X"01C9", X"00E4", X"044F", X"0517", X"02E9", X"0064", X"00DE", X"FDB8", X"FE37", X"FC69", X"FE30", X"01EF", X"0408", X"03CB", X"0207", X"00DE", X"0130", X"0041", X"FC2B", X"F7C4", X"FAE8", X"FCF7", X"000C", X"0267", X"00B1", X"FFB2", X"FD30", X"0220", X"020D", X"01AB", X"00BD", X"03DA", X"043D", X"01C9", X"0267", X"0165", X"004F", X"FF7C", X"0182", X"02FB", X"0478", X"02F1", X"030E", X"FFB0", X"015F", X"005D", X"FC82", X"FA8A", X"FADD", X"FF27", X"FFFC", X"016C", X"FEC6", X"FE89", X"FD4D", X"FCD8", X"02F8", X"0197", X"0011", X"017B", X"01FC", X"03E7", X"0656", X"05FD", X"0417", X"0313", X"0035", X"00FE", X"0196", X"007E", X"FFA6", X"FE08", X"021E", X"FCD3", X"F8C5", X"FABD", X"FE83", X"006D", X"0059", X"003E", X"00B5", X"FD75", X"FC89", X"FB01", X"FEEF", X"0008", X"FD08", X"FF3A", X"FFE1", X"02C7", X"0505", X"0747", X"038E", X"03C0", X"00D4", X"FF5D", X"0019", X"FEE0", X"FE42", X"FD32", X"FDBF", X"FF8F", X"F99E", X"FC2E", X"FF74", X"FF18", X"FF36", X"FF2A", X"04B7", X"0467", X"FEB2", X"FD01", X"FF35", X"FF22", X"FF78", X"00B1", X"FF79", X"0277", X"01B2", X"0460", X"03F2", X"03C8", X"032F", X"00C5", X"FFF5", X"FDFD", X"FDF9", X"FC21", X"FB6A", X"FE3F", X"FE17", X"FEBF", X"FC88", X"009C", X"FFAB", X"00C0", X"0018", X"05B7", X"03B6", X"FD8C", X"0160", X"01DB", X"02A9", X"055E", X"0532", X"0543", X"06B6", X"05F0", X"06CF", X"044A", X"0352", X"004C", X"FE96", X"FE9C", X"FD96", X"FC34", X"FCAD", X"FF93", X"FEB6", X"FB01", X"FCB1", X"0027", X"FE4D", X"00CC", X"0064", X"00CA", X"FE22", X"FDAC", X"008C", X"FFF5", X"0176", X"01F9", X"0269", X"0240", X"0250", X"00B0", X"FFF2", X"002E", X"0171", X"00E1", X"FE31", X"FFC7", X"FC4C", X"FF03", X"02C9", X"0376", X"0406", X"FD61", X"FD49", X"0095", X"FF72", X"FF56", X"00FE", X"FEEE", X"FFE7", X"FEE8", X"FDDC", X"FC0A", X"FBD0", X"FA61", X"FBF2", X"FF03", X"FE0F", X"FDC7", X"FD1F", X"FC17", X"FC30", X"FC4D", X"FACB", X"FB90", X"FF01", X"FF30", X"FED5", X"FE33", X"023F", X"FF57", X"004A", X"002A", X"FFBF", X"FEDF", X"FF25", X"008B", X"FF8A", X"FDB5", X"FDA2", X"FD9B", X"FD4B", X"FCC2", X"FF8A", X"003C", X"FFC7", X"FCCB", X"FD1E", X"FD6C", X"FA9A", X"FABD", X"F9CF", X"FA43", X"FBB5", X"F98C", X"FBD7", X"FE77", X"0052", X"FFB1", X"FFE1", X"FFF5"),
--        (X"0106", X"FE75", X"FF26", X"0010", X"0114", X"FFE6", X"0071", X"0093", X"FF69", X"FFD7", X"0016", X"001B", X"FFAE", X"FE84", X"FF92", X"0209", X"FF6F", X"FFA6", X"FF9D", X"0008", X"00B6", X"002A", X"FF89", X"FFB7", X"FF55", X"000B", X"FF9B", X"000A", X"0096", X"00B1", X"006A", X"FF03", X"00E1", X"00A8", X"FC54", X"FB46", X"FBB4", X"FCF6", X"FB05", X"FAFF", X"F850", X"FB27", X"00A8", X"0256", X"023A", X"FE5A", X"FB56", X"FBA0", X"FC43", X"FC20", X"FD40", X"003A", X"0095", X"FFF8", X"0049", X"FF85", X"FFC5", X"0060", X"0066", X"FF58", X"FEE6", X"FF44", X"FD60", X"FAA6", X"FB16", X"FF10", X"FACF", X"FE1E", X"FFCB", X"FF48", X"0030", X"02B0", X"03FB", X"02E8", X"0097", X"FC73", X"F997", X"F801", X"FA09", X"FB52", X"0059", X"0142", X"FF84", X"FF76", X"00DA", X"FF5A", X"0320", X"0169", X"FC3E", X"FF71", X"00FB", X"0000", X"0267", X"0345", X"037F", X"03BD", X"033E", X"058F", X"05B7", X"04F0", X"051B", X"02D2", X"FFF2", X"FE03", X"FB16", X"F8FA", X"F526", X"F4D7", X"F9A4", X"FF2F", X"FE4B", X"FF08", X"FF68", X"0041", X"03C4", X"01D6", X"0025", X"02B2", X"03FB", X"0374", X"0172", X"01EF", X"0129", X"0067", X"FEF1", X"012E", X"0136", X"01F6", X"0350", X"0090", X"FFF0", X"0101", X"FEE4", X"FB09", X"F9AB", X"F62D", X"F944", X"F9FA", X"FB9C", X"FDFF", X"012E", X"00B3", X"0269", X"0237", X"01BA", X"054D", X"02F8", X"01CC", X"FF60", X"0138", X"01E1", X"FE21", X"FE7E", X"FE88", X"FFF5", X"013C", X"0270", X"FF3D", X"0070", X"0093", X"FFD0", X"FE90", X"FDE2", X"FB1A", X"FAEF", X"F67B", X"FB63", X"FCC0", X"FFE6", X"025D", X"041E", X"071A", X"064D", X"0540", X"02F4", X"FFE0", X"FF48", X"0099", X"01AB", X"FFD6", X"FFF8", X"FFD9", X"0165", X"0139", X"0053", X"0081", X"0235", X"0072", X"0016", X"FED2", X"FCD0", X"FA7D", X"F82C", X"F3B5", X"FC4A", X"FEC2", X"00D4", X"0386", X"049E", X"0733", X"07E4", X"0416", X"01CE", X"00E7", X"00C2", X"02BB", X"03E8", X"0351", X"00BA", X"00B6", X"008C", X"0088", X"00AF", X"01F9", X"0325", X"01F4", X"012A", X"00F6", X"FE1D", X"FA23", X"F310", X"F38B", X"FDBE", X"FD16", X"FE24", X"0474", X"06D1", X"0812", X"0915", X"039D", X"043E", X"0420", X"059C", X"0387", X"0658", X"05D3", X"03FF", X"0149", X"00B6", X"0253", X"01D7", X"02E4", X"0318", X"015C", X"0212", X"004F", X"FF4C", X"F97B", X"F21B", X"F5C4", X"FBBD", X"0033", X"002C", X"03B0", X"084B", X"0893", X"065C", X"0625", X"0517", X"0561", X"048A", X"0533", X"0314", X"FFE8", X"FBA2", X"F960", X"FE8C", X"0392", X"0439", X"0213", X"0134", X"FEED", X"FFD9", X"FEE3", X"FFFA", X"FC2E", X"F38B", X"F64C", X"FC37", X"003B", X"015B", X"02EA", X"0745", X"069A", X"0127", X"0180", X"0009", X"FF68", X"FFFF", X"FDFE", X"F982", X"F691", X"F12A", X"F224", X"FB95", X"007D", X"0262", X"03D5", X"0129", X"FF8D", X"FF87", X"FF64", X"FC7E", X"FD40", X"F67A", X"FE5E", X"FE3E", X"029D", X"0289", X"01E7", X"05BA", X"019E", X"FB7E", X"F858", X"F617", X"F55C", X"F2A7", X"F1BB", X"F0DD", X"F112", X"F28A", X"F2EF", X"FBF8", X"00D8", X"0035", X"0110", X"00AB", X"0015", X"FFCC", X"FE18", X"FC24", X"FD72", X"FA4B", X"00E6", X"FEB6", X"FF36", X"0167", X"0171", X"0164", X"FC07", X"F4CB", X"EF72", X"EEF4", X"EBF4", X"EDDE", X"EE07", X"F4C5", X"F778", X"F8BE", X"FA23", X"FDB9", X"005C", X"0047", X"FDBC", X"FE36", X"FE0D", X"FC47", X"F9DC", X"FA90", X"F980", X"FFA8", X"07FD", X"0598", X"0307", X"0001", X"FF35", X"0192", X"FA52", X"F2D1", X"EB55", X"ECB2", X"EE94", X"F313", X"F910", X"FCE2", X"FFAC", X"FE1D", X"00ED", X"00CC", X"FEA1", X"FE85", X"FE84", X"FF50", X"FE62", X"FCD9", X"FDA6", X"FBEE", X"FC0B", X"011F", X"09F6", X"0BCF", X"02D7", X"0091", X"FEF0", X"028B", X"FA5F", X"F780", X"F229", X"F6B1", X"FBDF", X"FF12", X"023E", X"027A", X"0199", X"01D1", X"0474", X"03E5", X"00D8", X"FEBA", X"FEB7", X"00A1", X"006E", X"FF81", X"0051", X"FF4B", X"FFC1", X"027E", X"0873", X"0770", X"02AD", X"FF43", X"011E", X"0274", X"FEE4", X"FD7C", X"FED0", X"014F", X"017B", X"0209", X"03F2", X"02DE", X"02E0", X"01DC", X"02C2", X"02F0", X"0118", X"FEAE", X"FE87", X"0030", X"FF3F", X"FDEA", X"02B2", X"00B0", X"024F", X"0421", X"06A7", X"0B50", X"042A", X"0168", X"00AB", X"044D", X"03CA", X"037A", X"0348", X"0551", X"04E2", X"0238", X"019E", X"FFD6", X"01B3", X"0184", X"0619", X"02CF", X"FFE5", X"FF50", X"0169", X"FFBE", X"0132", X"001E", X"02C7", X"0258", X"038C", X"0724", X"09BD", X"0BA7", X"0354", X"012B", X"0066", X"0643", X"07FD", X"080B", X"03AA", X"028B", X"02A3", X"FF52", X"FFC8", X"FEF3", X"FE60", X"0049", X"025C", X"0195", X"FE84", X"FE88", X"005D", X"01C0", X"00DB", X"FFA0", X"011D", X"0208", X"0262", X"0444", X"0922", X"094F", X"035D", X"0192", X"019E", X"0342", X"092C", X"06EF", X"058A", X"0335", X"0032", X"FFB1", X"0027", X"FE60", X"FE1C", X"002F", X"027B", X"004F", X"FF46", X"0080", X"01C3", X"0169", X"01C1", X"0019", X"0174", X"02CA", X"0358", X"058A", X"07DC", X"073D", X"02FC", X"FF6E", X"FD51", X"FF84", X"0648", X"0668", X"0211", X"012E", X"02F3", X"FFC9", X"FFA1", X"FDBE", X"FD72", X"FF07", X"01B7", X"0073", X"FEDB", X"FFDA", X"00B2", X"FF84", X"FEC1", X"FFAC", X"011B", X"FF36", X"0071", X"00C1", X"0771", X"07A8", X"01DB", X"0011", X"FF1C", X"00FE", X"06F7", X"0778", X"035E", X"036C", X"0154", X"00BB", X"0151", X"FFE3", X"0055", X"FE46", X"FEE2", X"FE3D", X"FDD6", X"FE17", X"FFCF", X"0031", X"00F3", X"FF3D", X"FE72", X"FEF1", X"FFE9", X"0279", X"065E", X"0675", X"0057", X"FF52", X"012E", X"04FF", X"0546", X"0495", X"0320", X"03EF", X"01B8", X"00BA", X"FFE0", X"004E", X"FFA7", X"FC3F", X"FCE5", X"FE36", X"FE74", X"FEBC", X"FE37", X"FEBD", X"00B7", X"FEAE", X"FE4B", X"FE88", X"0013", X"002E", X"027A", X"01CF", X"FFA1", X"FFBA", X"013A", X"05DE", X"03E9", X"0544", X"058D", X"05EB", X"0292", X"FFF4", X"FEC2", X"FDB0", X"FD96", X"FBAB", X"FE30", X"FCBD", X"0018", X"FEFD", X"FFAE", X"01EE", X"026E", X"FFFA", X"00C4", X"008E", X"001D", X"FFC4", X"FF09", X"FDFD", X"006B", X"FF7A", X"FF75", X"044A", X"00C9", X"04CC", X"06A6", X"0491", X"0152", X"FEFE", X"FE53", X"FE57", X"FFA5", X"FD5B", X"FE8F", X"FE55", X"FEAB", X"FF1A", X"FE08", X"0227", X"FFFF", X"FE06", X"FD06", X"00CF", X"FE72", X"FF8E", X"FF87", X"00E5", X"0026", X"008B", X"FF9E", X"03B4", X"01EB", X"06A7", X"0470", X"0536", X"03FA", X"0115", X"FFA1", X"009F", X"00EB", X"01BD", X"FF5D", X"00A9", X"FDCC", X"FC7D", X"FE38", X"FBFA", X"FA59", X"FDCC", X"FDAF", X"FEB9", X"FE58", X"03AD", X"022B", X"0283", X"FFAC", X"005A", X"0086", X"FE75", X"FE13", X"0301", X"006C", X"FF22", X"026A", X"0577", X"05D9", X"04FB", X"0495", X"0589", X"0350", X"00B1", X"0177", X"FF27", X"FCF5", X"FAFC", X"F8F0", X"F903", X"F89F", X"F9CB", X"FACD", X"FECA", X"01BF", X"01A6", X"FFD7", X"FFE8", X"0031", X"FFAB", X"FFE2", X"FB0B", X"FD30", X"FDEA", X"007E", X"02F4", X"032B", X"03C9", X"01E3", X"02AC", X"0095", X"0110", X"0396", X"01C5", X"0133", X"FFCA", X"FF86", X"FDDB", X"FA99", X"FBE6", X"FD98", X"0186", X"0034", X"0076", X"FF8F", X"006A", X"0021", X"017C", X"00E2", X"01E2", X"0147", X"0175", X"0391", X"0239", X"025A", X"0428", X"0589", X"0642", X"07AA", X"055D", X"07D0", X"0654", X"058D", X"0291", X"016D", X"FEAA", X"FE6E", X"FDFA", X"00FF", X"FEFF", X"FFF0", X"FF65", X"002F"),
--        (X"0127", X"003E", X"0062", X"FFD3", X"01CE", X"FEBF", X"FFDF", X"008C", X"0020", X"FF34", X"FF2E", X"000C", X"00D4", X"0000", X"FF14", X"FF9A", X"0116", X"FF02", X"013F", X"017F", X"0010", X"FED4", X"FFE2", X"00CB", X"00BA", X"007E", X"FE49", X"FEBD", X"002D", X"004D", X"0006", X"FF5E", X"000A", X"FFB5", X"02D3", X"028D", X"02F2", X"03AD", X"0324", X"0410", X"0421", X"03B0", X"FD47", X"FD93", X"FE42", X"0071", X"0133", X"0122", X"01BB", X"00E5", X"00A4", X"01D2", X"FF9F", X"FF36", X"FEA6", X"FE63", X"003F", X"0033", X"FFB0", X"FFE7", X"000D", X"018C", X"038F", X"03C3", X"03D8", X"01F7", X"0401", X"0245", X"03B4", X"FEC9", X"004C", X"FE17", X"013E", X"00C5", X"0387", X"04FA", X"03EA", X"0411", X"01AF", X"020F", X"0090", X"FEF6", X"FF93", X"0023", X"00AD", X"01BA", X"FF3C", X"00EE", X"024E", X"FCB6", X"FDCF", X"FDBC", X"FF10", X"FE0B", X"FD8F", X"FAE6", X"FA14", X"FB93", X"FCEB", X"FF14", X"FF84", X"0152", X"04CD", X"07A8", X"07AD", X"078D", X"04D5", X"00E5", X"02EF", X"0125", X"023C", X"00DF", X"007D", X"0036", X"FCEC", X"FD77", X"FAB5", X"FBE7", X"FD06", X"FD37", X"F89D", X"F9A9", X"FC57", X"FC94", X"FBF3", X"F9B8", X"FCD5", X"FE62", X"FFDE", X"0310", X"0131", X"01BE", X"0352", X"04BF", X"0569", X"06AF", X"0517", X"FFC8", X"FD86", X"0110", X"00AF", X"FE59", X"0025", X"FC3B", X"F98D", X"F8F3", X"FBF4", X"FC98", X"FDAF", X"FF5D", X"FF4E", X"FE89", X"FCC0", X"FCF0", X"FD57", X"FB8E", X"FF1C", X"FFF3", X"017D", X"FF46", X"0275", X"0436", X"0589", X"05F8", X"0317", X"FFEA", X"0105", X"01DC", X"0011", X"FD93", X"01AD", X"FC63", X"F987", X"FD2D", X"FEF9", X"0032", X"FF7D", X"FED5", X"FE8B", X"FDAA", X"FE0A", X"FCA6", X"FE45", X"FE46", X"FD35", X"FFFF", X"002F", X"0268", X"0121", X"03F7", X"068D", X"05D9", X"0579", X"FDCA", X"0107", X"014D", X"019D", X"FD56", X"029D", X"FCCB", X"F80F", X"FD49", X"FF79", X"003F", X"011C", X"009F", X"0090", X"013F", X"FE28", X"FCDA", X"FE56", X"FCF7", X"FF4E", X"0193", X"01EE", X"025A", X"0094", X"041E", X"08B0", X"08AE", X"06D3", X"0579", X"02CB", X"0217", X"02DF", X"03F2", X"05D3", X"FD75", X"F6B0", X"FD1F", X"009C", X"00C8", X"0336", X"0348", X"0205", X"0201", X"0152", X"FCDC", X"FB5B", X"FC5C", X"FDB1", X"FDFF", X"FDFF", X"FE94", X"FF3F", X"02E1", X"059D", X"0BA2", X"0ABA", X"0664", X"006B", X"FEFC", X"01A4", X"0445", X"0776", X"FD7F", X"F9F4", X"FDE5", X"0198", X"0131", X"01D0", X"03B2", X"031A", X"0333", X"0393", X"005E", X"FC74", X"F7C4", X"F9DA", X"FA7E", X"FE6E", X"FBEE", X"FE82", X"032E", X"0778", X"0BE0", X"0D56", X"085F", X"0236", X"02EA", X"0192", X"02E7", X"0528", X"FD75", X"FFCC", X"0232", X"0144", X"0420", X"053A", X"0616", X"053E", X"028F", X"030B", X"0202", X"FC67", X"FB44", X"FB76", X"FA95", X"FAB0", X"F8A6", X"FE00", X"03E2", X"080A", X"0C6E", X"0DDA", X"079B", X"01F6", X"0024", X"0057", X"05E6", X"04D4", X"00CA", X"0220", X"031E", X"0362", X"04A5", X"0534", X"040F", X"0253", X"0028", X"027F", X"FF36", X"FB75", X"FB49", X"FBE1", X"FBFB", X"FA17", X"F9CA", X"FD41", X"0507", X"0AD0", X"0CE3", X"0A8E", X"0716", X"FFB2", X"FE49", X"01AD", X"0338", X"0785", X"01F0", X"0191", X"0196", X"032E", X"02E2", X"013B", X"FE50", X"0064", X"000B", X"0367", X"FD4C", X"F9B4", X"FA93", X"FAFE", X"FA76", X"FA2B", X"FE60", X"0128", X"096C", X"0B1B", X"0A5E", X"04D6", X"001F", X"FEFB", X"FF4F", X"FEAC", X"0137", X"04A3", X"0237", X"04A6", X"0415", X"01BF", X"0004", X"FE04", X"FD9B", X"01BD", X"03A1", X"021E", X"FABA", X"FA54", X"F9DA", X"F96E", X"FB98", X"FEBA", X"0496", X"090D", X"0CF4", X"0AF5", X"0852", X"0554", X"010F", X"FD2A", X"FDBC", X"015C", X"FF95", X"03A4", X"FF9D", X"04F1", X"0728", X"015F", X"01C7", X"FFB7", X"00A7", X"038C", X"046E", X"00DF", X"FAC4", X"FACA", X"FA06", X"FCB2", X"FF24", X"0303", X"06F2", X"0ACF", X"0A4C", X"09EB", X"05BE", X"05BA", X"FFFA", X"FB76", X"00BF", X"0184", X"FD51", X"FF7C", X"FD29", X"02FA", X"077D", X"03DC", X"008A", X"FF90", X"0116", X"04DF", X"04D2", X"00F9", X"FC44", X"F970", X"FC9E", X"0118", X"04DF", X"0679", X"06C4", X"07D0", X"05D7", X"059D", X"0450", X"02EB", X"FEAB", X"FD78", X"FDE6", X"FF0A", X"FB9C", X"FA0F", X"FC07", X"0118", X"05E5", X"02C9", X"015F", X"0060", X"FDA0", X"0180", X"02CC", X"FD90", X"FB99", X"FD72", X"00F0", X"047C", X"04B3", X"0464", X"0609", X"065A", X"03AD", X"021E", X"00DC", X"FF81", X"FF0D", X"FBAB", X"FD68", X"0061", X"FD1A", X"FAA7", X"F9D7", X"FF18", X"04D5", X"0748", X"015F", X"FF36", X"FF14", X"0088", X"008A", X"FEDC", X"FD3A", X"019A", X"0440", X"03E8", X"053B", X"063C", X"01FC", X"02EA", X"00CD", X"FE97", X"FE73", X"FF2E", X"FD7F", X"FBB7", X"FC46", X"003F", X"FFE8", X"FD19", X"F992", X"0180", X"0641", X"0596", X"0270", X"FFB6", X"FF50", X"002A", X"0296", X"00FF", X"0232", X"0466", X"01EB", X"025D", X"0302", X"0058", X"017D", X"FF0E", X"FD91", X"FC3E", X"FCCB", X"FFC6", X"FDB7", X"FDF5", X"FC72", X"FE5B", X"0303", X"0265", X"FADB", X"0186", X"0288", X"01EE", X"02F7", X"0202", X"FF70", X"00E9", X"04D0", X"0481", X"0209", X"02D0", X"0265", X"FF5D", X"FE50", X"FEE9", X"FC92", X"FD9B", X"FD62", X"FBDC", X"FE37", X"FFCF", X"FD20", X"FC02", X"FDE4", X"0148", X"0165", X"02AA", X"FDB9", X"FEE9", X"0197", X"0096", X"FEE8", X"FEE0", X"00FB", X"023E", X"0546", X"03B8", X"0188", X"0151", X"0098", X"FFD3", X"FD50", X"FBA5", X"FDC7", X"FB0F", X"FB44", X"FE29", X"FDCF", X"FE3C", X"FEF0", X"FCF3", X"FE86", X"0015", X"FF6D", X"FEB1", X"FD1B", X"FFFE", X"025D", X"FF5E", X"FF35", X"0087", X"0127", X"0183", X"04F1", X"0334", X"01FB", X"00AA", X"FFD9", X"FE52", X"FD2A", X"FD9B", X"FB09", X"FD56", X"FEE3", X"005D", X"FED8", X"00DE", X"FDA8", X"0305", X"FFBD", X"FFDE", X"FF3C", X"FC6F", X"FC39", X"006E", X"FF76", X"FF80", X"FF4B", X"0065", X"00C2", X"0157", X"01E8", X"0177", X"0182", X"00A4", X"0119", X"0188", X"FF08", X"FD6B", X"FDB3", X"FE77", X"FDFC", X"FF69", X"013F", X"00E0", X"FEC2", X"024E", X"FF62", X"FF5A", X"005F", X"FBD0", X"FC93", X"FD88", X"011A", X"00EE", X"FF4C", X"0114", X"0132", X"01A4", X"0125", X"FF43", X"FFF0", X"0265", X"0150", X"0026", X"FF2B", X"FC51", X"FDDE", X"FDF8", X"00AD", X"00B9", X"0088", X"FDDC", X"FF88", X"021C", X"FF7C", X"0150", X"00A8", X"FCFF", X"FCD0", X"F9FE", X"FE95", X"FFFA", X"0045", X"024F", X"020F", X"0119", X"00BE", X"0061", X"022F", X"024A", X"0140", X"0182", X"00A7", X"FFC4", X"FD2F", X"FDE3", X"FF1F", X"01A4", X"0107", X"001A", X"FDA2", X"FFC3", X"00CA", X"00E8", X"0084", X"FEBC", X"0220", X"00E9", X"FFB6", X"FDAC", X"FDF8", X"FE4C", X"0144", X"001D", X"01F2", X"001D", X"FFA4", X"0181", X"01E7", X"01E4", X"00EF", X"FFCF", X"FF77", X"FA2F", X"FD05", X"0154", X"03B0", X"025D", X"002E", X"0108", X"FEE4", X"003E", X"003E", X"FFE6", X"FFEE", X"FFBC", X"0238", X"03B0", X"FFFD", X"00E7", X"FEA9", X"FF2A", X"FECC", X"FF90", X"009D", X"FCEF", X"00BE", X"FC49", X"FAA4", X"FD8A", X"FEBA", X"FB86", X"FC3D", X"FCE2", X"FAF5", X"FFB8", X"00E5", X"FF8A", X"FF97", X"00A4", X"FEF3", X"003C", X"FFC1", X"FF58", X"013C", X"007D", X"0082", X"00A8", X"0114", X"0070", X"FE6A", X"009C", X"03BF", X"FA4D", X"FCDE", X"028B", X"03E0", X"007C", X"01B1", X"0103", X"FD07", X"FD54", X"011A", X"012A", X"00C6", X"00F6", X"012E"),
--        (X"0292", X"0021", X"FDCE", X"0071", X"FFDA", X"FEFF", X"FEB2", X"FFCC", X"FF28", X"FED4", X"FF05", X"FFCE", X"00D3", X"FF68", X"0044", X"FF87", X"0130", X"FF34", X"FF0D", X"01C2", X"00AA", X"00F0", X"FFFD", X"015A", X"FF0C", X"FFDF", X"FF0C", X"FF37", X"00D0", X"FFAB", X"FF4D", X"010D", X"FF49", X"0014", X"007A", X"01DA", X"00D6", X"0090", X"0066", X"04BB", X"03F6", X"0292", X"FE0B", X"FD3F", X"02DC", X"0400", X"FFF9", X"FFEE", X"FFA0", X"FFD5", X"00DB", X"FF89", X"FEA0", X"FF83", X"FFC6", X"FF10", X"FE1A", X"FFF8", X"0119", X"FF30", X"FF5F", X"FF4E", X"FF20", X"0366", X"02EA", X"016A", X"0370", X"0662", X"0525", X"00C5", X"0009", X"FBFA", X"FF1E", X"0156", X"00B1", X"00FD", X"0223", X"04E7", X"0190", X"0231", X"042A", X"0273", X"FF00", X"FF8F", X"008B", X"FEC1", X"FE07", X"FE3C", X"FDF3", X"0357", X"02B1", X"04E8", X"0453", X"02DD", X"03D1", X"03CE", X"046C", X"0279", X"0283", X"FE4F", X"FF57", X"0077", X"00F1", X"01A7", X"FFE3", X"FD41", X"FEB4", X"0012", X"0196", X"01D7", X"0089", X"0086", X"00A2", X"0124", X"FDCF", X"FD94", X"002D", X"04A9", X"057E", X"0551", X"065A", X"079B", X"05CF", X"050B", X"0413", X"0393", X"0037", X"FF6F", X"01AC", X"00AA", X"0038", X"FC16", X"FE1F", X"FBB0", X"FD56", X"FAC8", X"FB05", X"FF6A", X"01A5", X"025E", X"0088", X"0027", X"FF73", X"FEAD", X"01CC", X"FF69", X"FF91", X"0232", X"03FD", X"021C", X"043C", X"047F", X"0541", X"0460", X"01C5", X"01AB", X"02F7", X"04BC", X"04BD", X"01B5", X"013E", X"FE96", X"FD31", X"F9D0", X"FB4E", X"00F4", X"FFAA", X"0269", X"007F", X"006C", X"FF73", X"FE9A", X"FF91", X"FDD4", X"FD72", X"00C1", X"0169", X"0216", X"005F", X"00AE", X"01C3", X"0346", X"0254", X"0213", X"03A0", X"01FD", X"017F", X"00D2", X"0176", X"FF0E", X"FD82", X"FE59", X"FCE9", X"FF61", X"FDFB", X"FCF5", X"FF0B", X"0041", X"FE7B", X"FB3B", X"01B1", X"FF2D", X"FF7D", X"FF90", X"0203", X"FEAB", X"FFC5", X"FF33", X"FF74", X"0037", X"0044", X"015E", X"00C4", X"FE26", X"FD43", X"FE25", X"FD81", X"FE12", X"FE3B", X"FEAA", X"FE54", X"FF98", X"FF18", X"FC00", X"027E", X"FD62", X"FBC9", X"FC0D", X"FF45", X"FEAF", X"FC4A", X"FE0F", X"FD6C", X"FF18", X"00A1", X"FDD7", X"FDB8", X"FDBA", X"FC1D", X"FCB2", X"FDDE", X"FD42", X"FAC3", X"FC3A", X"FC89", X"FDF3", X"FDED", X"FED8", X"FDE9", X"FD06", X"0069", X"FFCE", X"FEC4", X"FC30", X"FD51", X"FC86", X"FE65", X"FE9D", X"FE51", X"FF60", X"008F", X"01DF", X"0278", X"019D", X"FE1C", X"FD48", X"FBEE", X"FC5C", X"FBB9", X"FAF2", X"FC94", X"FC11", X"FE5B", X"FDE6", X"FD38", X"FF18", X"F909", X"F773", X"FCD7", X"FBBE", X"FE52", X"FC6C", X"FA0D", X"FEBB", X"FCA8", X"FDA0", X"0162", X"00A3", X"0176", X"0219", X"0383", X"0195", X"FE6F", X"F9AA", X"FA67", X"F9AF", X"F803", X"FB67", X"FBB5", X"FE7D", X"FF4E", X"FE68", X"FFF3", X"FEBB", X"F828", X"F3B1", X"F969", X"FD40", X"FFB1", X"FB09", X"F9D8", X"FCAE", X"FD96", X"FF64", X"0285", X"0169", X"037D", X"04D5", X"0710", X"0550", X"FDF3", X"F7D3", X"F950", X"F981", X"F959", X"FE3F", X"00BE", X"02E9", X"0452", X"00F3", X"0303", X"0377", X"FEFF", X"F4F6", X"FB6D", X"FC16", X"FE41", X"FB2C", X"F8A4", X"FB31", X"FBED", X"FFA8", X"00D2", X"FDEC", X"FE89", X"02AC", X"07EF", X"0896", X"04DA", X"FF30", X"FDD7", X"FD69", X"005A", X"02E8", X"04B3", X"05FC", X"07AB", X"0942", X"0ADE", X"0943", X"0CBE", X"FC44", X"FC8A", X"FF4E", X"FE8F", X"FE38", X"F9DB", X"FF39", X"FB31", X"FE5B", X"FD23", X"FE88", X"FF6E", X"0244", X"07B7", X"0704", X"0758", X"06A1", X"031E", X"011E", X"036B", X"04B6", X"049D", X"06A7", X"0638", X"096F", X"0BB5", X"06F7", X"071E", X"026D", X"03CB", X"0229", X"FE68", X"FEBF", X"FAC9", X"FF0C", X"FDD7", X"FCCB", X"FEE0", X"010A", X"01BF", X"0315", X"04C2", X"043F", X"0717", X"067A", X"03AA", X"01AA", X"0194", X"030B", X"FE7A", X"FFFF", X"018D", X"050B", X"03FB", X"0304", X"0521", X"031C", X"03BD", X"010A", X"FD96", X"0128", X"FC29", X"FEA6", X"FF88", X"0034", X"FFC2", X"0020", X"0022", X"0324", X"03E6", X"03ED", X"05BC", X"037A", X"004D", X"FF84", X"017C", X"FEBE", X"FCD8", X"0028", X"0100", X"0116", X"0130", X"02D5", X"05AB", X"06A3", X"0451", X"01D1", X"FFD0", X"003E", X"01EF", X"000B", X"02AA", X"030D", X"FEA4", X"FFD9", X"0247", X"03BE", X"0463", X"0671", X"05D0", X"0117", X"FEF1", X"FE00", X"025D", X"FF3E", X"009D", X"01CC", X"0181", X"0155", X"03D4", X"06AD", X"0780", X"08CB", X"01F9", X"01B0", X"008A", X"00A1", X"02E4", X"0297", X"01A8", X"00C7", X"0188", X"00C1", X"022C", X"03CC", X"04D4", X"05F2", X"01D1", X"FF67", X"FBE7", X"FD53", X"0160", X"01E2", X"026A", X"02EA", X"0097", X"02D9", X"0373", X"0322", X"0398", X"066D", X"0058", X"0302", X"FF8A", X"FFC0", X"FD4E", X"023A", X"02D8", X"0122", X"007B", X"FFEE", X"0071", X"003E", X"0260", X"0356", X"FF8B", X"FD80", X"FB87", X"FDB2", X"FFE4", X"018F", X"0343", X"01F9", X"007B", X"03B4", X"0606", X"0488", X"05B9", X"0469", X"FE20", X"FE1E", X"FFCB", X"FC1F", X"FDDF", X"059C", X"03ED", X"0506", X"0217", X"FFC1", X"FF02", X"FEC0", X"013F", X"008E", X"FE30", X"FC9C", X"FAF3", X"FE28", X"019E", X"0261", X"03A6", X"01A0", X"0219", X"05BC", X"064A", X"0602", X"00F4", X"FFBE", X"FED1", X"FDF6", X"002D", X"01A6", X"018C", X"0440", X"061B", X"03C6", X"0240", X"00F6", X"FD1F", X"FDDC", X"FF9A", X"FF6B", X"FDA5", X"FCD3", X"FC5B", X"FFBF", X"FFE1", X"0120", X"02F6", X"02BE", X"05DA", X"056D", X"0650", X"074C", X"045E", X"01DE", X"FDCD", X"FF0C", X"FF4A", X"00CD", X"0640", X"03F0", X"0234", X"00AE", X"0010", X"FEB9", X"FBFB", X"FE63", X"FE03", X"FFD8", X"0033", X"FF01", X"FCCF", X"FEA3", X"FFD9", X"000D", X"03C5", X"0493", X"046D", X"0445", X"0911", X"09B4", X"04EC", X"01E9", X"00C6", X"FF27", X"FFF2", X"00A7", X"05B8", X"04F1", X"FFD9", X"FDCB", X"FF2E", X"FD91", X"FEC1", X"FF33", X"FFC0", X"00F9", X"033C", X"0435", X"FEE3", X"FE82", X"005D", X"0086", X"0313", X"03A3", X"04FB", X"0661", X"0A01", X"078B", X"02CB", X"0198", X"FCC1", X"0102", X"FFB5", X"0015", X"0328", X"076F", X"FEE5", X"FD6D", X"FC7C", X"FF00", X"02BC", X"FFF6", X"00A4", X"0293", X"0243", X"04A3", X"027E", X"002E", X"00DE", X"015D", X"0313", X"0776", X"068B", X"0721", X"09FC", X"095A", X"04F7", X"037F", X"FEC9", X"FF63", X"0156", X"015D", X"021A", X"0006", X"008D", X"FC28", X"FD8A", X"FEC1", X"FFCB", X"FFF7", X"003F", X"0159", X"0186", X"02FC", X"030D", X"02AB", X"0694", X"0255", X"0526", X"04FC", X"0374", X"0581", X"0530", X"0617", X"0376", X"0035", X"000A", X"FEF1", X"FF88", X"0051", X"01F3", X"FD40", X"FE73", X"FEC4", X"FF67", X"0015", X"FDE5", X"FDA1", X"FEFF", X"FDC1", X"FBC0", X"FEE6", X"00C0", X"FFB7", X"021D", X"FF95", X"FEFB", X"FEFF", X"0012", X"0001", X"FFD6", X"03C3", X"FFAD", X"FFCD", X"0196", X"0095", X"00F0", X"00E1", X"FF84", X"006D", X"020B", X"0199", X"029D", X"03A5", X"01BC", X"01DB", X"FFFE", X"FFBE", X"003C", X"FF8A", X"00B3", X"FF0D", X"FDF4", X"FE10", X"FA74", X"F942", X"FE6A", X"FF74", X"FEC1", X"FF85", X"FF98", X"0034", X"001D", X"006E", X"FE7C", X"FF19", X"FF8D", X"FEBC", X"00A7", X"FF47", X"0207", X"01E8", X"FEB8", X"FFEC", X"FE37", X"0068", X"FFB6", X"FAC6", X"FE28", X"FECF", X"FBD3", X"F96B", X"FC1E", X"FC26", X"FEF3", X"FFAD", X"FF82", X"FB78", X"0148", X"00A7", X"FF47", X"0111"),
--        (X"FFD8", X"00BA", X"FF44", X"FF90", X"006B", X"00D1", X"0057", X"0051", X"FE91", X"FFC4", X"FE08", X"FFBA", X"FE11", X"FE06", X"006C", X"FE53", X"FEAC", X"FEDA", X"FFA7", X"FFDD", X"FED9", X"FF46", X"FEB1", X"0097", X"0032", X"0015", X"FF2E", X"FFE8", X"003C", X"0009", X"0046", X"00A6", X"FE70", X"FDFE", X"FC12", X"FB65", X"FB6F", X"FB49", X"FB7B", X"FA1A", X"F878", X"F9BE", X"FBA4", X"F9FC", X"FA32", X"FACF", X"FA57", X"FA48", X"FA01", X"FBC6", X"FDA6", X"FC33", X"0013", X"FF8C", X"00D1", X"005E", X"004D", X"FFA5", X"0011", X"FD9C", X"FE55", X"FE62", X"F901", X"F922", X"F64B", X"F548", X"F3A0", X"F278", X"F348", X"F43C", X"F0FF", X"F3BB", X"FA02", X"FD68", X"FD5E", X"FE2F", X"FC46", X"FD62", X"FEB4", X"FAEC", X"FD3E", X"FF0D", X"015B", X"000C", X"008F", X"00A6", X"FF3B", X"FEBF", X"0140", X"FC2B", X"FB59", X"F90F", X"F86A", X"F95D", X"F8FB", X"F669", X"F7A9", X"F699", X"F72B", X"FC66", X"FBA4", X"FF5A", X"0241", X"0086", X"0321", X"0423", X"FF72", X"FB3E", X"FE32", X"FCEE", X"FE70", X"0049", X"00F1", X"005E", X"FFB9", X"0288", X"FECF", X"0069", X"0130", X"FFC3", X"FE84", X"FE6F", X"FE54", X"FE64", X"FDBE", X"FC27", X"FD61", X"FEF1", X"FEFE", X"0128", X"0215", X"0098", X"FDF1", X"02B2", X"02E9", X"0290", X"044B", X"01FD", X"FF01", X"FDF7", X"0001", X"0018", X"FCF9", X"0223", X"FD35", X"031A", X"0345", X"0265", X"037D", X"01CD", X"02BC", X"0116", X"FF1E", X"FC67", X"FD56", X"FD95", X"FE62", X"FEE4", X"FE4D", X"FF4C", X"FE0B", X"FF42", X"02F7", X"037E", X"01B8", X"0226", X"03E8", X"FFDF", X"00BB", X"01F6", X"0040", X"0093", X"FE61", X"02F4", X"03E2", X"03E6", X"047F", X"04E6", X"0693", X"0444", X"0156", X"FF3B", X"00BA", X"FDD6", X"00B1", X"FF06", X"FEB4", X"FED6", X"FFB4", X"FFD7", X"FE7E", X"00A0", X"03CF", X"02E7", X"04B3", X"FF21", X"0197", X"03F4", X"FF1D", X"03E8", X"FE99", X"0328", X"03F4", X"04C1", X"0612", X"04BC", X"0317", X"047F", X"0391", X"0314", X"02AB", X"FFDF", X"00A9", X"000C", X"FFE8", X"0130", X"02D6", X"0006", X"0055", X"00F2", X"0242", X"0591", X"02A8", X"007C", X"FD5B", X"FFBE", X"FFDC", X"0255", X"FE54", X"02DF", X"02D8", X"03E0", X"0363", X"02AE", X"0407", X"022F", X"0160", X"00B7", X"00D1", X"00E7", X"FEBE", X"0028", X"0108", X"0084", X"044F", X"017D", X"02AF", X"0343", X"0538", X"08A2", X"030D", X"FFA7", X"00AF", X"030F", X"0065", X"0060", X"005B", X"02C7", X"025F", X"02C6", X"00C8", X"00D8", X"00C4", X"0079", X"00E4", X"FF54", X"FED3", X"0061", X"FF2B", X"00AB", X"0213", X"FEEA", X"0103", X"0295", X"023E", X"012F", X"09EF", X"0A70", X"05D5", X"0179", X"FF9A", X"0082", X"FF52", X"01EB", X"004B", X"0246", X"018D", X"01CE", X"0169", X"009B", X"00B3", X"0123", X"0220", X"0092", X"FE87", X"0064", X"0303", X"006E", X"0133", X"FFF7", X"0017", X"FEAF", X"FE20", X"FC84", X"040D", X"0C62", X"069C", X"0100", X"00A5", X"FE9B", X"038E", X"025F", X"0130", X"008E", X"0223", X"0081", X"0277", X"FFD1", X"00FB", X"0322", X"041A", X"00D7", X"FD79", X"01EA", X"038F", X"03FE", X"01D0", X"FE4F", X"F9FF", X"F9C5", X"F8C4", X"F743", X"F9D3", X"038D", X"0539", X"0193", X"FFAC", X"FF78", X"009F", X"02B7", X"00ED", X"0212", X"0144", X"0207", X"02ED", X"01ED", X"0347", X"04E2", X"01EE", X"FEE1", X"FE49", X"FFCE", X"0351", X"0392", X"015E", X"FE1C", X"FAB3", X"F7BA", X"FA0C", X"F4CD", X"F2FE", X"FC9A", X"034C", X"0024", X"FEB6", X"FFFE", X"0170", X"013C", X"0306", X"0305", X"018D", X"02F4", X"0292", X"0390", X"049C", X"034C", X"007E", X"FE6E", X"FD21", X"FD79", X"020B", X"04C6", X"0181", X"FE3F", X"FDF9", X"FD0A", X"FC0B", X"F8D6", X"F796", X"F96F", X"FBD5", X"FC46", X"00B9", X"02ED", X"0267", X"01D1", X"0374", X"003E", X"FF25", X"013C", X"0240", X"0120", X"0161", X"FF06", X"0079", X"FD75", X"FDF5", X"01C8", X"0557", X"03A6", X"0089", X"FE3B", X"FE3D", X"006E", X"00EB", X"0028", X"FC46", X"F8BD", X"FC6B", X"FDE0", X"FE8A", X"00FB", X"0083", X"020E", X"FF0B", X"FBCA", X"FBBB", X"FBA7", X"FF58", X"FF0C", X"0072", X"0089", X"FF60", X"FEF1", X"FDE1", X"01F8", X"0485", X"0562", X"0096", X"0026", X"FF04", X"02AC", X"01DD", X"0359", X"FE72", X"F8FB", X"0022", X"FC85", X"FE54", X"0193", X"0210", X"FE71", X"FBEA", X"FC67", X"F900", X"F8C0", X"FA79", X"FA3C", X"FAC5", X"FE11", X"0033", X"0148", X"01F4", X"035A", X"04AB", X"02B8", X"018E", X"0274", X"0196", X"0247", X"030A", X"02EE", X"0033", X"F7C9", X"FDCD", X"FB33", X"FFFD", X"0243", X"03E7", X"FFE1", X"FF5D", X"FC1E", X"FD7E", X"F9CC", X"F7BC", X"FA3D", X"F796", X"F9CF", X"FB89", X"FF93", X"02DC", X"0604", X"043D", X"036E", X"0348", X"0032", X"00D8", X"01F8", X"00FE", X"0153", X"FE84", X"F9BC", X"FE11", X"FBD7", X"0037", X"0218", X"04FA", X"0460", X"0100", X"FF26", X"FF97", X"FDEA", X"FB08", X"F917", X"F757", X"F991", X"F9C9", X"0161", X"0467", X"060E", X"0325", X"030D", X"FF93", X"0103", X"0114", X"FFF9", X"FE88", X"FD7E", X"FC60", X"F88C", X"02C3", X"FEBA", X"FF60", X"FDB4", X"070C", X"064B", X"0238", X"0120", X"0149", X"FE96", X"FEC1", X"FC2E", X"F8A7", X"F972", X"FA14", X"FEDA", X"02E5", X"0060", X"0053", X"FEB9", X"005A", X"FF90", X"00DF", X"FDBE", X"FBB9", X"FDC7", X"FF96", X"FAFE", X"FC38", X"FD27", X"FF96", X"FF62", X"049F", X"071F", X"0163", X"005E", X"FF98", X"FB1B", X"FEB6", X"FD9D", X"FAE3", X"FACA", X"FACD", X"FF06", X"FF35", X"FD36", X"00DB", X"FF55", X"FF8B", X"00A9", X"FF6C", X"FDEF", X"FCE0", X"FDD1", X"FEF8", X"007B", X"FDD1", X"FF46", X"0093", X"0085", X"001F", X"0381", X"0084", X"FF99", X"FD1D", X"FD46", X"00BE", X"FCA9", X"FDB7", X"FD62", X"FE50", X"FEF1", X"FD25", X"FF13", X"FF8D", X"FEE9", X"FF7A", X"010F", X"FF27", X"008B", X"FF1D", X"FF78", X"FFA9", X"0048", X"FDF4", X"0031", X"FF81", X"FF95", X"0179", X"015F", X"0122", X"FB2B", X"FC51", X"FC3C", X"FE1C", X"FD23", X"FEAC", X"FEEE", X"FE98", X"FDDA", X"FDD6", X"FF01", X"FE71", X"0095", X"01A1", X"01F0", X"016E", X"00EA", X"FFE4", X"0023", X"00B0", X"00E4", X"003B", X"0104", X"00A3", X"016E", X"014A", X"069B", X"04E8", X"0418", X"014D", X"00FC", X"FE6F", X"FD0F", X"FFB3", X"01B6", X"FDB6", X"FC0D", X"FE08", X"FE66", X"FE79", X"FF3D", X"0083", X"039F", X"070A", X"055E", X"FFE3", X"0132", X"0153", X"0346", X"02D9", X"FFD9", X"0050", X"FFEB", X"017D", X"0733", X"0994", X"0A72", X"07D5", X"07B3", X"0220", X"00FB", X"0144", X"000C", X"FD31", X"FE0D", X"FED5", X"FF3D", X"FF85", X"01A9", X"03B3", X"0664", X"06C7", X"058E", X"04FE", X"05D3", X"0001", X"FDB2", X"FDCB", X"01CE", X"FF7D", X"FEE6", X"0172", X"0381", X"08D0", X"0A5A", X"0762", X"09A7", X"079E", X"06C9", X"05FB", X"0524", X"06A6", X"0704", X"05ED", X"088E", X"06A0", X"08D9", X"0877", X"0759", X"0580", X"06A9", X"0813", X"068D", X"045E", X"FCB6", X"FD4A", X"FF39", X"00D3", X"FF00", X"FF97", X"00FD", X"0210", X"0364", X"03EF", X"046E", X"0375", X"0538", X"0460", X"064C", X"04C1", X"0673", X"069F", X"067E", X"06BF", X"077C", X"0523", X"00F2", X"02D9", X"0604", X"045C", X"FFBE", X"FEE1", X"001B", X"FE68", X"FF6B", X"FF2C", X"FEA9", X"00FD", X"0027", X"00D9", X"01E4", X"FFEB", X"00DD", X"015A", X"00D6", X"02F6", X"02C2", X"01EC", X"0374", X"0378", X"03E4", X"02C8", X"FFF2", X"0081", X"FFF1", X"020A", X"04CF", X"0281", X"021D", X"FFEC", X"FF8F", X"FFF1", X"FFD8"),
--        (X"FF4C", X"008E", X"FFAB", X"FEFA", X"00DA", X"FFF4", X"FF60", X"FF01", X"FFA1", X"0047", X"FEE0", X"FF84", X"FEFF", X"0055", X"007A", X"FF2F", X"FEFF", X"01AD", X"FF98", X"FF1D", X"FF63", X"FE69", X"003B", X"0031", X"0059", X"00C4", X"FEEC", X"FFC7", X"FF7C", X"0031", X"FFCE", X"FF1D", X"FE26", X"FECA", X"FECB", X"001C", X"FEF4", X"0058", X"0084", X"FE5E", X"FDD6", X"FDD2", X"01B2", X"0210", X"FBEB", X"FC94", X"0129", X"0199", X"FFDB", X"00C6", X"FEFC", X"00B2", X"00ED", X"004E", X"FFF1", X"FFF0", X"0116", X"0061", X"01B4", X"FF4A", X"FEC0", X"00FC", X"FD5A", X"FE9A", X"FA08", X"FB2C", X"FD6C", X"0064", X"00F0", X"00B9", X"00A2", X"0589", X"05A8", X"0326", X"FE4A", X"FD9B", X"FF31", X"FDD7", X"FEFD", X"FEC6", X"FEE6", X"0037", X"FFE6", X"00BF", X"FF86", X"0124", X"01A4", X"00C9", X"FF0B", X"0242", X"021A", X"0041", X"0086", X"0060", X"004E", X"FF8A", X"0409", X"01EC", X"015C", X"0403", X"0395", X"00D8", X"007C", X"024B", X"0330", X"FE0A", X"FADE", X"F831", X"F9C5", X"FE6D", X"FE1D", X"0112", X"0005", X"0128", X"028A", X"03D7", X"0389", X"0416", X"024E", X"0251", X"0454", X"00DD", X"012D", X"0033", X"FFAA", X"00D9", X"FFDC", X"FEA9", X"FF36", X"FCAD", X"FF04", X"01A1", X"00BE", X"01E5", X"FFFC", X"FC7D", X"F83E", X"F870", X"FC18", X"FC94", X"FF65", X"FFD6", X"0147", X"0326", X"0528", X"0830", X"048D", X"0477", X"01FC", X"0172", X"FF92", X"FE11", X"FC74", X"FA0A", X"FBA0", X"FC81", X"FC3A", X"FB60", X"FC34", X"FF5B", X"0054", X"FE71", X"FD89", X"FCFF", X"FD7C", X"F501", X"FB47", X"FD8F", X"008D", X"015E", X"0143", X"0460", X"0650", X"0610", X"059A", X"0285", X"01BF", X"01A9", X"FFBD", X"FE9D", X"FDB4", X"FE93", X"FCFE", X"FD9B", X"FE5A", X"FD87", X"0062", X"0001", X"020D", X"022F", X"0058", X"FDE2", X"FB05", X"F438", X"F941", X"FF25", X"001F", X"01FE", X"FFD2", X"071F", X"0A7C", X"05C0", X"054D", X"03EF", X"0105", X"00A5", X"009E", X"FEC5", X"0057", X"FFBA", X"017B", X"0211", X"0209", X"01E1", X"0266", X"0251", X"04C7", X"0206", X"00B1", X"FD76", X"F957", X"F650", X"FB88", X"FD51", X"FCD7", X"00A5", X"02CF", X"05EA", X"0B51", X"07EE", X"0311", X"011C", X"FEF5", X"FEF2", X"FEBF", X"FDDC", X"FFD9", X"0203", X"0414", X"0666", X"03C4", X"032A", X"0282", X"0246", X"01D9", X"013C", X"02D6", X"FEA6", X"F887", X"F8DD", X"FC28", X"FDE1", X"009D", X"0161", X"04EB", X"046B", X"0702", X"055A", X"0170", X"FFB3", X"FD6F", X"FC22", X"FBA3", X"FBC5", X"FEB9", X"02CF", X"07DE", X"0819", X"051D", X"02EE", X"0291", X"0213", X"03D6", X"0349", X"03B7", X"FD96", X"F88A", X"F744", X"FBDC", X"00EB", X"00DB", X"0368", X"0344", X"050E", X"0169", X"FFBB", X"FEB8", X"FEAF", X"FBB4", X"FABF", X"FB3F", X"FBA3", X"FBC3", X"0578", X"08F2", X"0696", X"0548", X"043C", X"0315", X"0174", X"049C", X"0273", X"0354", X"FDB5", X"F766", X"FE09", X"FD1F", X"006D", X"0008", X"0455", X"0334", X"0583", X"0172", X"FEC1", X"FDB5", X"FCA6", X"FB74", X"FBA4", X"FC0E", X"FE15", X"00A2", X"05FE", X"0884", X"066F", X"059A", X"0493", X"0397", X"027D", X"0244", X"026C", X"00DC", X"FDF1", X"F56C", X"FB5B", X"FDF8", X"0159", X"0163", X"01AA", X"03AB", X"0310", X"01FF", X"FE3C", X"FD7F", X"FD81", X"FE2B", X"FDBD", X"FEDF", X"FE19", X"FFC3", X"0377", X"06DC", X"0593", X"03D5", X"031B", X"0241", X"FF95", X"FE4C", X"FC3E", X"FC77", X"FB21", X"F829", X"FE5F", X"FFB7", X"02EE", X"007C", X"00F9", X"02A8", X"024B", X"033E", X"FE5C", X"FEE3", X"FF1C", X"FE94", X"FD68", X"FD61", X"FCD6", X"FBAC", X"0249", X"04BB", X"027C", X"0291", X"0135", X"FEEF", X"00CC", X"FDA1", X"FD04", X"FA15", X"FC68", X"FC99", X"FF8D", X"FB6C", X"FC95", X"FE29", X"00DB", X"03A6", X"FEED", X"008E", X"00FB", X"FF44", X"FE58", X"FC72", X"FDC9", X"FBA4", X"FA5D", X"FD62", X"FFE1", X"0317", X"014E", X"009C", X"0023", X"01D4", X"01E2", X"FF57", X"002E", X"FFBC", X"00BE", X"FE6E", X"FC5A", X"F8B6", X"FDF8", X"FD14", X"01CB", X"01CC", X"FF57", X"0071", X"00BF", X"004C", X"FD72", X"FAEF", X"FAE0", X"FB68", X"FC5E", X"FCE5", X"FF03", X"0073", X"0228", X"FEAB", X"FF7D", X"0030", X"020D", X"01D8", X"0154", X"0390", X"0261", X"FE3C", X"F73B", X"FD0B", X"FD10", X"015D", X"02F9", X"0142", X"00ED", X"0320", X"0183", X"FFDF", X"FFB0", X"FBF3", X"FBD5", X"FCA1", X"FB80", X"FAE2", X"FE8A", X"01AB", X"008D", X"FF68", X"FFE4", X"01E3", X"014F", X"019A", X"01B7", X"0385", X"01DF", X"FDBF", X"F11B", X"FAD2", X"FC0B", X"016A", X"039A", X"0032", X"0355", X"0439", X"0144", X"FC5B", X"FC79", X"F9A4", X"FA3E", X"F81E", X"FA46", X"F9CA", X"FED5", X"017E", X"00D5", X"00A2", X"FF33", X"01B6", X"0157", X"0013", X"0273", X"02D4", X"0321", X"FB2E", X"F696", X"FED1", X"FB98", X"0288", X"0186", X"0254", X"03EC", X"04C0", X"0183", X"FE41", X"FB17", X"FAFF", X"FA72", X"F971", X"F97F", X"F9CF", X"FDC3", X"00E8", X"01D0", X"006A", X"01FE", X"00DC", X"015A", X"0127", X"022D", X"02CD", X"FD01", X"F424", X"F79A", X"0211", X"008D", X"0095", X"0211", X"0135", X"0537", X"05B7", X"0111", X"FF03", X"FD00", X"FD34", X"FDD9", X"FBB7", X"F98B", X"FBD1", X"0055", X"02DC", X"0126", X"0022", X"FFDA", X"0030", X"FFD8", X"FF9F", X"000A", X"FE60", X"F8CA", X"F6EB", X"FC26", X"FFA7", X"01B2", X"FFF7", X"FE6C", X"FDED", X"02E1", X"038C", X"00F7", X"0092", X"FF4D", X"FFCA", X"FEA2", X"FD95", X"FD3F", X"FD5F", X"FEF9", X"01C8", X"FF3E", X"021A", X"0144", X"FF9A", X"FDCE", X"FF85", X"FD71", X"FC14", X"F7F5", X"F7D2", X"FBFC", X"004B", X"011D", X"FEC0", X"FE4C", X"FF2A", X"0058", X"0299", X"FFE3", X"01A4", X"FFD9", X"01A9", X"FFF9", X"FF3D", X"FF0D", X"FD73", X"FEC1", X"001E", X"015F", X"0047", X"006F", X"FFDD", X"FF0A", X"FCA1", X"FCD8", X"F9A3", X"F438", X"F75A", X"FCDC", X"FE84", X"008D", X"0168", X"FFF4", X"003F", X"FE84", X"00D8", X"03ED", X"0341", X"0293", X"025B", X"00A0", X"0003", X"FD1C", X"FBF2", X"FB05", X"FE6A", X"01C9", X"FFA6", X"0179", X"0271", X"014F", X"FE7D", X"F93A", X"F7DD", X"F4DF", X"F704", X"FA9F", X"026F", X"FF83", X"0179", X"0081", X"00A0", X"02C4", X"03E6", X"0708", X"083F", X"0755", X"02BF", X"026A", X"0107", X"FF93", X"FFFF", X"FDC8", X"FDC2", X"FFA0", X"FF36", X"FF1E", X"0111", X"FD29", X"F8AA", X"F73E", X"F6F5", X"F659", X"F9EA", X"FBF3", X"03C7", X"00B9", X"FE4B", X"0089", X"FFAC", X"0422", X"0684", X"08BD", X"0A18", X"0A02", X"07FD", X"064D", X"030A", X"FF87", X"FF8E", X"019D", X"FFDB", X"FED2", X"FE33", X"FD1F", X"FC56", X"F8A9", X"FA4F", X"FAFB", X"FB2B", X"F6D4", X"FB39", X"FDFD", X"0191", X"FFCC", X"FE11", X"FF98", X"FE5D", X"0142", X"03B5", X"06F2", X"0630", X"0785", X"0976", X"0930", X"061F", X"0896", X"0663", X"0479", X"03F3", X"01A6", X"0136", X"013A", X"01C8", X"001C", X"FD5E", X"FF4A", X"00F3", X"FC33", X"FFD1", X"FF02", X"0060", X"FFBA", X"0071", X"FF67", X"0038", X"0026", X"FF2D", X"00FE", X"02B0", X"0379", X"0320", X"049C", X"0288", X"00F1", X"FF42", X"009A", X"039E", X"02BF", X"0409", X"0600", X"0509", X"049C", X"019C", X"01CB", X"024F", X"0206", X"00E2", X"0071", X"FF09", X"0072", X"005E", X"0014", X"016B", X"008C", X"009C", X"0014", X"0013", X"FF78", X"0013", X"031E", X"014C", X"01B9", X"00FE", X"03EF", X"012D", X"0353", X"0371", X"0334", X"020C", X"FFF9", X"FF10", X"FF70", X"00C1", X"03C6", X"005C", X"00BE", X"0078", X"006C"),
--        (X"00FD", X"016D", X"FEF8", X"0061", X"0125", X"FFB4", X"0125", X"013B", X"FDEA", X"00E0", X"FF9C", X"0094", X"FF96", X"FFD4", X"0041", X"0160", X"0012", X"00ED", X"0137", X"FF70", X"FFC5", X"0026", X"FF8D", X"0051", X"014D", X"0010", X"0028", X"FF70", X"0066", X"0125", X"00B6", X"004E", X"001E", X"FF25", X"FDEF", X"FD59", X"FC53", X"FF82", X"FF9E", X"FF5F", X"FD00", X"FB3E", X"FDC9", X"FE40", X"FEEB", X"FE8E", X"FCF0", X"FD87", X"FCAC", X"FF9C", X"FF37", X"FF72", X"014C", X"FEA3", X"FF92", X"FF09", X"0120", X"FFD6", X"FF93", X"FF12", X"FEEC", X"000C", X"FE98", X"FD57", X"0088", X"0316", X"0325", X"025E", X"0098", X"FE7A", X"FE17", X"FA3A", X"F99D", X"F716", X"F8FD", X"F861", X"F910", X"F99E", X"F8F9", X"FB14", X"FD6F", X"FF11", X"0076", X"001D", X"0023", X"0055", X"FDBE", X"FD7B", X"FD3D", X"FF88", X"FFD2", X"01C0", X"0421", X"0557", X"05D2", X"0348", X"01D6", X"018C", X"0164", X"FD1C", X"FAE6", X"FAD9", X"F8D5", X"F745", X"F675", X"F852", X"FA0D", X"FCCF", X"FD8B", X"014D", X"FFEE", X"0012", X"FFF0", X"FF51", X"FE2B", X"FC05", X"FDB4", X"FD5B", X"FE5B", X"FF82", X"013F", X"0472", X"0463", X"0263", X"0239", X"010D", X"FFE7", X"FD1B", X"FF92", X"FF58", X"FFA6", X"FF62", X"007D", X"FF1E", X"FFAD", X"FE3C", X"FD30", X"FDF0", X"FFED", X"0088", X"FFDB", X"008F", X"FEB2", X"FFED", X"FEA6", X"FDBF", X"FE7A", X"0036", X"02C4", X"01BE", X"017B", X"0092", X"012A", X"FEF4", X"FFC9", X"FE5F", X"00A0", X"01B0", X"00A0", X"0140", X"0253", X"0400", X"001A", X"FECA", X"FEB1", X"FE07", X"FD65", X"FF92", X"FFF6", X"FFAA", X"FF21", X"01D4", X"000C", X"FE99", X"00E2", X"02B6", X"0331", X"01BB", X"017D", X"00E6", X"FEBF", X"FE58", X"FDC1", X"FF19", X"FE97", X"FF47", X"FCDF", X"0081", X"0149", X"02E6", X"0226", X"FFC3", X"FE36", X"FD35", X"FDAA", X"FF59", X"0273", X"FE0C", X"03BD", X"0283", X"0085", X"00C7", X"0097", X"0157", X"0151", X"01EA", X"0300", X"0034", X"FFEA", X"FE98", X"FB5E", X"FD00", X"FDAB", X"FDEA", X"001C", X"FFAA", X"005B", X"FE8C", X"01C9", X"0239", X"FF5B", X"FE74", X"0103", X"FE38", X"0032", X"0159", X"04E5", X"039A", X"0160", X"0071", X"01C3", X"0135", X"0027", X"0163", X"017E", X"007B", X"016B", X"FE4F", X"FCA9", X"FC94", X"FE46", X"0070", X"01E4", X"0137", X"008B", X"FFEB", X"0116", X"02D3", X"FEA5", X"FB30", X"FE47", X"FE77", X"011B", X"03E5", X"02FC", X"02B0", X"0069", X"013B", X"FF2C", X"0026", X"FF21", X"FFC6", X"014B", X"00D0", X"00C1", X"0035", X"FF26", X"0043", X"04D1", X"0576", X"0466", X"0367", X"02B8", X"0310", X"0106", X"FF7F", X"FAFC", X"F956", X"FE11", X"FE49", X"00AD", X"0350", X"0302", X"FF65", X"01F4", X"0364", X"0132", X"FF60", X"FDA2", X"0110", X"0122", X"00F1", X"0079", X"FEC6", X"FF3D", X"0236", X"0618", X"04EB", X"043D", X"042D", X"0490", X"0293", X"0377", X"02A9", X"FA65", X"F85E", X"F87A", X"FE0C", X"0031", X"042B", X"0553", X"00EC", X"0278", X"0239", X"0339", X"0034", X"FFD9", X"01A2", X"002C", X"FFC4", X"FEB5", X"FD5D", X"FDF7", X"009F", X"0233", X"02EC", X"02CD", X"0345", X"0391", X"05C8", X"06D6", X"028C", X"FC11", X"FB0B", X"F9A2", X"FC6D", X"0156", X"02E5", X"05F9", X"0472", X"0316", X"02F3", X"024E", X"FE91", X"FF17", X"FF77", X"FEED", X"FEE4", X"FDCE", X"FBF9", X"FCB5", X"FF4D", X"FFEE", X"0123", X"FEFB", X"02EA", X"031E", X"0741", X"0794", X"0701", X"077A", X"01E5", X"FF3B", X"0200", X"FEA9", X"02C3", X"0419", X"0621", X"025B", X"0121", X"0396", X"FFA0", X"FE64", X"FF3C", X"FDCE", X"FFDE", X"0033", X"FD85", X"FE5B", X"FE65", X"FEA8", X"0094", X"FFAA", X"00B2", X"0281", X"04D5", X"078C", X"0B7A", X"0942", X"0764", X"0551", X"013D", X"FE62", X"FFD4", X"01A5", X"0606", X"03D2", X"06CC", X"0699", X"01CD", X"FED2", X"FB14", X"FCB1", X"FF36", X"FEDB", X"FD0B", X"FE10", X"FCFA", X"FF26", X"014D", X"01F6", X"0119", X"0112", X"FFA9", X"03FD", X"08B2", X"0A16", X"05F8", X"044C", X"011E", X"0023", X"FCD9", X"FDEA", X"0297", X"07FA", X"0A18", X"0902", X"0AB6", X"0382", X"FC43", X"F9BF", X"F947", X"FAB6", X"FBCA", X"FFC8", X"FF83", X"0143", X"0240", X"0239", X"0052", X"FFBE", X"FC74", X"FC4F", X"0662", X"09C9", X"060C", X"03AD", X"02A2", X"00CB", X"FC87", X"FDEA", X"005D", X"077C", X"0CF1", X"0F3F", X"0FCC", X"0EAA", X"079B", X"001A", X"FBC7", X"FCA6", X"FEE0", X"015D", X"0223", X"0051", X"02BC", X"0167", X"00EF", X"FF35", X"FCC6", X"FBC6", X"036C", X"09B5", X"08AF", X"055D", X"01D3", X"00E3", X"FF2A", X"001E", X"FDDB", X"0163", X"07CE", X"0D2A", X"0F14", X"12B4", X"12C1", X"0D3D", X"0852", X"0759", X"06E2", X"0278", X"0214", X"028A", X"0222", X"FF9C", X"FE68", X"FE54", X"FC02", X"FF0F", X"02D1", X"0A77", X"084E", X"0480", X"0255", X"00FC", X"FF7F", X"FF67", X"FA43", X"FE30", X"0341", X"04FE", X"0AD8", X"0FCC", X"1296", X"126B", X"11AE", X"0F5E", X"0977", X"0405", X"00BC", X"00C9", X"FED8", X"FEF7", X"FD61", X"FF0F", X"FD6D", X"FF68", X"03FE", X"08F0", X"0632", X"023E", X"FEE9", X"002C", X"01E9", X"FF37", X"FAC5", X"FC55", X"FDA3", X"FD87", X"0271", X"0523", X"0951", X"0B5F", X"0999", X"08BC", X"05EC", X"00E5", X"FF76", X"FE97", X"FFFE", X"FEF0", X"FEE5", X"FECD", X"FD86", X"FED2", X"0207", X"045C", X"0339", X"0227", X"000D", X"FF63", X"00AE", X"FD30", X"FA59", X"FC02", X"FD00", X"FB0A", X"FC49", X"FB1C", X"FDFB", X"003E", X"0000", X"0265", X"FF54", X"FF90", X"FF41", X"FF8D", X"FEB4", X"FE8B", X"00BE", X"FE60", X"FF95", X"FF5D", X"FE3B", X"02AD", X"02F5", X"FF83", X"FF9F", X"FECC", X"FEC7", X"FFE0", X"FAE9", X"FAEB", X"FB9C", X"FB97", X"FCAC", X"FB50", X"FC2F", X"FCA8", X"FDA0", X"FE3A", X"FEA0", X"FFDD", X"004A", X"FF61", X"FEA9", X"FF8D", X"FE6F", X"FDAC", X"FF0A", X"FF90", X"00BD", X"025C", X"0328", X"01DA", X"00BC", X"FE61", X"FE7C", X"FF1E", X"FDFD", X"FA2C", X"FD57", X"FE9B", X"FEDC", X"FDC3", X"FBFC", X"FD5E", X"FD85", X"FF12", X"FFF7", X"0095", X"0134", X"FF71", X"FED5", X"FF5D", X"FE79", X"FC66", X"FFF8", X"00F8", X"FE1F", X"03B1", X"054D", X"FC8A", X"00AB", X"FFA2", X"FFCB", X"FD25", X"F8AB", X"F969", X"FBCD", X"FDA6", X"FFC8", X"FDC9", X"FCE2", X"FB9C", X"FDBD", X"FDD6", X"FF43", X"002D", X"0035", X"FF53", X"0025", X"FFC1", X"FFC6", X"FFDD", X"01A0", X"03D9", X"01B3", X"00F4", X"02AC", X"FD31", X"FF57", X"FEFD", X"FF9D", X"002C", X"F932", X"F7C9", X"F9FE", X"FA7D", X"FB2D", X"FBD7", X"FBDD", X"FB66", X"FE20", X"FED2", X"FF1D", X"0013", X"0287", X"0023", X"FEFE", X"00AB", X"0236", X"00C5", X"008D", X"FE7F", X"FE31", X"02BB", X"0144", X"FF4B", X"FF89", X"0019", X"FFC7", X"FED9", X"013B", X"FF6B", X"FA73", X"F966", X"FA44", X"F89B", X"F9CA", X"FA5A", X"FCB3", X"FCB9", X"FC26", X"FE86", X"0074", X"FE0A", X"0067", X"0255", X"003F", X"FEB1", X"FDFD", X"FC7D", X"FB95", X"FDBC", X"FD1D", X"00E8", X"FF7F", X"00D0", X"014B", X"0019", X"FFB5", X"FAB2", X"FAD3", X"FBA6", X"FD01", X"FE0C", X"FC2E", X"FBD9", X"FB7D", X"FC62", X"FE44", X"FB14", X"FF42", X"FEAE", X"FF99", X"FEC6", X"025E", X"FDAB", X"FF5D", X"FFDF", X"FE38", X"001F", X"FF98", X"0140", X"FFE1", X"00C3", X"FFCE", X"FFDA", X"FEDD", X"00BC", X"FFDD", X"0152", X"0184", X"01E6", X"0126", X"FF2E", X"FF69", X"FE55", X"024A", X"FC83", X"FF19", X"00FD", X"01E8", X"0126", X"011E", X"0477", X"02A1", X"035F", X"001F", X"FFC0", X"0085", X"FE89", X"001D"),
--        (X"FF8F", X"000F", X"FF44", X"FFC5", X"FFF2", X"FE5F", X"FFC9", X"FF8B", X"0038", X"FFB0", X"FFF2", X"0074", X"02BD", X"010D", X"002F", X"FFED", X"FF98", X"00F8", X"FFF5", X"FFC3", X"FECE", X"FFB2", X"FFBB", X"006A", X"0005", X"002A", X"FF90", X"006A", X"FFA4", X"00C3", X"FF99", X"001F", X"002F", X"00AE", X"03A3", X"0323", X"032E", X"04F7", X"065D", X"058C", X"0731", X"0869", X"0232", X"0717", X"02EC", X"055D", X"060A", X"05C5", X"057E", X"0304", X"0264", X"01E6", X"FF77", X"FF00", X"0075", X"0086", X"FFA7", X"FF96", X"FF2B", X"0308", X"0374", X"0295", X"053D", X"06FA", X"0604", X"023B", X"0197", X"047B", X"0828", X"08DE", X"0968", X"063F", X"043F", X"03FA", X"04AD", X"08BF", X"05F3", X"05BA", X"06E1", X"04BE", X"FECC", X"FFE0", X"0109", X"FDD8", X"0098", X"001A", X"015B", X"01EB", X"0442", X"040C", X"0299", X"00AC", X"009C", X"0136", X"FFA6", X"016B", X"0405", X"0595", X"0311", X"0286", X"03F8", X"0158", X"03E2", X"062A", X"03BF", X"044E", X"0289", X"02FD", X"0199", X"FE5F", X"02CC", X"0082", X"00A4", X"00C8", X"0109", X"02C0", X"0474", X"0029", X"FF2A", X"FFB4", X"FF4D", X"FEF6", X"00D1", X"FEA4", X"FFA0", X"FDDB", X"FF30", X"0218", X"026B", X"01EC", X"02C5", X"01CC", X"FDE5", X"FF7E", X"0336", X"02C2", X"024C", X"0168", X"FE26", X"006F", X"0109", X"FFAF", X"FEEF", X"FFA1", X"FDD1", X"FF8E", X"0156", X"FF10", X"FE3E", X"FEAE", X"001F", X"FD42", X"FE82", X"FFB9", X"FE5C", X"0058", X"00C7", X"0287", X"0123", X"FFF3", X"FEDE", X"FCB4", X"025C", X"01AE", X"0065", X"FE7F", X"027A", X"011D", X"0039", X"FF24", X"0160", X"FD6E", X"FE95", X"0142", X"FFD5", X"FE31", X"FE4E", X"FD7F", X"FE3A", X"007D", X"FE1B", X"0145", X"004B", X"0009", X"0023", X"020A", X"00E8", X"FF8E", X"FD99", X"0031", X"002F", X"023D", X"0365", X"031F", X"024E", X"FFB1", X"FF20", X"0054", X"FD2D", X"FD6E", X"FE34", X"FE99", X"FE0B", X"FD13", X"FE4A", X"FE71", X"FF3B", X"0058", X"005D", X"FF1F", X"01F9", X"0183", X"02A0", X"03EC", X"0132", X"FC93", X"FD7D", X"FD40", X"FE8D", X"0088", X"01D6", X"038D", X"00BF", X"0112", X"027D", X"FF2D", X"FAA1", X"FB48", X"FC8A", X"FB1E", X"FAF5", X"FBCB", X"FCFA", X"FECA", X"005A", X"FEC6", X"0095", X"FF00", X"00EB", X"0544", X"044B", X"0260", X"FDCC", X"FC7C", X"FD43", X"FD10", X"FD9E", X"022B", X"0527", X"0304", X"FF78", X"FF94", X"FF73", X"0022", X"FBFD", X"FD49", X"FC06", X"FADB", X"FCB1", X"FD93", X"FD5C", X"FC41", X"FDC9", X"FE8C", X"FFAA", X"0153", X"0641", X"0626", X"0293", X"FD64", X"FAE9", X"F87E", X"FB8A", X"FAF7", X"FC8C", X"0079", X"0608", X"075B", X"0244", X"0399", X"00EC", X"FFEA", X"FE45", X"FBAF", X"FC29", X"FAD6", X"FD09", X"FD07", X"FCCC", X"FD9F", X"FEF0", X"FFC5", X"030E", X"079F", X"0A70", X"0605", X"FF42", X"F9C0", X"F840", X"F9E3", X"FAFC", X"FCA7", X"FB8E", X"02F3", X"078F", X"0874", X"052B", X"FEAC", X"00EF", X"FE2A", X"FE04", X"FBC1", X"FD62", X"FCAF", X"FFDD", X"003B", X"FDFD", X"FFA6", X"0173", X"02CC", X"05C2", X"08BD", X"073E", X"FF05", X"F971", X"F894", X"FA32", X"FB6F", X"FAFB", X"FC13", X"FD0B", X"01FB", X"048F", X"04F3", X"01F6", X"FF2C", X"FF26", X"FC36", X"FEE8", X"FC85", X"FED8", X"0100", X"03F6", X"026C", X"0210", X"02B5", X"054F", X"06B4", X"082B", X"059B", X"00D7", X"FBF8", X"F615", X"F85E", X"F9E7", X"F895", X"F8F2", X"F849", X"FC71", X"FF7C", X"013A", X"FCF7", X"FBFC", X"FD7D", X"0059", X"000D", X"0058", X"026B", X"01AE", X"05CE", X"0617", X"05EF", X"03DB", X"0387", X"05EC", X"0430", X"031E", X"FFAD", X"FD80", X"F7CE", X"F9A6", X"F9C6", X"FA53", X"FAA9", X"F922", X"FBEA", X"FEE2", X"0375", X"01FC", X"FA1E", X"F75F", X"FE95", X"0415", X"0003", X"0117", X"FDCA", X"01B0", X"063C", X"0421", X"044A", X"046A", X"04B2", X"0643", X"FFF3", X"FE07", X"FCD8", X"FCEB", X"FB8E", X"FB28", X"F9DF", X"FC1E", X"FC4D", X"FCD5", X"FFEE", X"0288", X"064A", X"0446", X"FA4C", X"F951", X"FDE1", X"02F5", X"016B", X"009D", X"FA1D", X"FE6B", X"0324", X"0147", X"00CE", X"0308", X"0398", X"027E", X"002D", X"FCF3", X"FC86", X"FC27", X"FB53", X"FBA4", X"FBAC", X"FED7", X"0061", X"0128", X"0039", X"02B4", X"05FF", X"0449", X"FBE0", X"F891", X"FC59", X"FF3E", X"00EA", X"0007", X"FC69", X"FFAE", X"FDD6", X"FD89", X"FE43", X"0092", X"01BF", X"FF54", X"FE69", X"FB5B", X"F96B", X"FCA9", X"FB28", X"FB17", X"FA9E", X"FE4B", X"0025", X"012F", X"0205", X"02D8", X"0460", X"010B", X"FAF8", X"F893", X"FEDA", X"00E0", X"0140", X"FF08", X"FECA", X"FC37", X"FE9F", X"FDE1", X"FDA2", X"FE57", X"FF74", X"00B4", X"FCE0", X"F91F", X"F9B7", X"FAD5", X"FA40", X"FBDD", X"FCE1", X"FFA1", X"01D8", X"0283", X"02DC", X"04D7", X"0383", X"FD51", X"FBB2", X"FAFB", X"0192", X"FF16", X"0102", X"0114", X"0065", X"FCD1", X"FE74", X"000A", X"000C", X"01DB", X"0157", X"0091", X"FCCE", X"FA7F", X"FC42", X"FD87", X"FDB6", X"FEF3", X"0046", X"00D8", X"0123", X"02F0", X"0378", X"03D4", X"01FE", X"FEE1", X"FB38", X"FC64", X"FE1D", X"FFEB", X"03DC", X"02E4", X"0286", X"FE81", X"FD6D", X"FFE2", X"FE1D", X"FF2A", X"0026", X"02A0", X"0370", X"0201", X"0225", X"00BD", X"01E1", X"02AC", X"02B4", X"034D", X"0136", X"03B3", X"0314", X"0191", X"FF4D", X"002A", X"FCEF", X"FC8E", X"0079", X"FFF5", X"03AC", X"0109", X"0128", X"FE4F", X"FF00", X"FF72", X"FB92", X"FF14", X"01D8", X"0388", X"0318", X"0418", X"0371", X"03D5", X"0358", X"0451", X"0537", X"02C9", X"02FC", X"0258", X"0172", X"026E", X"01D2", X"FF40", X"0046", X"008B", X"FFA7", X"0135", X"00B4", X"0207", X"FEA4", X"FE8E", X"FE9C", X"FDD6", X"FC6E", X"FDEE", X"0063", X"0112", X"023F", X"02E7", X"0173", X"01F6", X"0281", X"02BC", X"02B4", X"02F4", X"016E", X"02FB", X"0069", X"0115", X"010C", X"FE1D", X"FF6C", X"0178", X"FF9C", X"0103", X"0192", X"01CB", X"004A", X"FE2D", X"FE7E", X"FF12", X"FDF1", X"FE94", X"FFB6", X"FF44", X"00C1", X"0082", X"0130", X"00C0", X"0179", X"030D", X"0360", X"0453", X"04C3", X"0173", X"014F", X"0067", X"FFB4", X"FE1E", X"FE11", X"0487", X"FFB9", X"0053", X"0076", X"02EC", X"04BD", X"0250", X"0073", X"FEE5", X"FE4D", X"FF84", X"0260", X"04C8", X"02B4", X"0330", X"00B7", X"027A", X"0188", X"027E", X"033C", X"016E", X"0187", X"0199", X"FD22", X"FE4C", X"FCAC", X"FD89", X"FEE7", X"0516", X"003E", X"0338", X"FFCD", X"00E2", X"0377", X"020B", X"037B", X"007D", X"023A", X"00B0", X"0221", X"00D1", X"FF8D", X"0126", X"0221", X"024F", X"0186", X"FFCF", X"024E", X"FFE2", X"0090", X"FD22", X"FF08", X"0019", X"0092", X"FECE", X"FEB0", X"00C9", X"00A6", X"FFC0", X"005F", X"0078", X"01C3", X"038E", X"00E5", X"FC6C", X"0086", X"FF3F", X"021B", X"FDA4", X"FEEF", X"FED6", X"FFCE", X"FBFD", X"FDEB", X"FF27", X"FFAD", X"FE4C", X"FF19", X"FE3B", X"0057", X"02E1", X"0305", X"032F", X"FFD7", X"FF91", X"0065", X"00BD", X"00F9", X"FF9F", X"FE33", X"FE29", X"FCFB", X"FA67", X"FA0B", X"F807", X"FB19", X"FAAF", X"004F", X"FF74", X"FF19", X"FD03", X"FE3C", X"FCCE", X"FCFF", X"FED9", X"FF7B", X"000E", X"FE33", X"009B", X"FED9", X"FD2A", X"FF40", X"FFC0", X"0113", X"FF58", X"FF8D", X"FF71", X"00E1", X"FFFC", X"FF01", X"FF39", X"FF86", X"FE51", X"FD0D", X"001C", X"00A0", X"0019", X"FED4", X"FC02", X"FB4D", X"FB4B", X"FBB7", X"FD82", X"FD90", X"00B6", X"0139", X"FCCF", X"FF5A", X"FDF0", X"0083", X"FF50", X"FED3"),
--        (X"0007", X"FF84", X"000E", X"FFFC", X"00BB", X"FF94", X"008C", X"017D", X"00EE", X"0167", X"FFC0", X"0056", X"0079", X"0194", X"0063", X"0146", X"0058", X"0046", X"00CA", X"0059", X"FFA2", X"FEF3", X"0140", X"01AE", X"0047", X"FF6F", X"FF39", X"FF71", X"FF7E", X"0121", X"0048", X"00FA", X"0007", X"FFDC", X"030A", X"01EB", X"036F", X"0471", X"03FF", X"04B5", X"0409", X"0216", X"00D0", X"041B", X"04F2", X"0501", X"0462", X"05B9", X"05B4", X"032E", X"0474", X"02DF", X"0131", X"0142", X"FF03", X"FFA0", X"FF0F", X"0133", X"FF32", X"014E", X"046E", X"002F", X"0217", X"04C6", X"0508", X"0821", X"07AD", X"09FB", X"06A6", X"0712", X"07A4", X"099A", X"080B", X"0692", X"0771", X"0688", X"0693", X"0918", X"059D", X"062A", X"0480", X"0192", X"0170", X"FFAA", X"0002", X"0103", X"FF85", X"0169", X"025B", X"0521", X"0488", X"08ED", X"0999", X"05C7", X"0865", X"06C9", X"0755", X"0A24", X"0A84", X"0A76", X"0A1B", X"0912", X"083E", X"06B8", X"0892", X"07F7", X"07FD", X"080E", X"06B6", X"FF52", X"FDD9", X"FE36", X"0090", X"FF69", X"FD76", X"00C2", X"FED7", X"FEF6", X"017E", X"045D", X"0469", X"02F8", X"03B0", X"0363", X"03E4", X"01DD", X"0427", X"0355", X"0482", X"04B3", X"04BC", X"02BC", X"039C", X"0437", X"0133", X"FDB4", X"FE37", X"FB85", X"FF78", X"0195", X"FF67", X"000F", X"0202", X"FFC2", X"FF6A", X"FCC3", X"0136", X"00E4", X"025A", X"013F", X"043B", X"046D", X"03F5", X"0397", X"0263", X"01C0", X"048E", X"05D3", X"078A", X"04B6", X"0154", X"0051", X"FDE8", X"FB35", X"FBD2", X"FF16", X"FF91", X"015A", X"FE19", X"009B", X"00D0", X"02DE", X"FD79", X"FC3E", X"0008", X"01ED", X"055F", X"03B0", X"03BB", X"0310", X"04CB", X"050C", X"0471", X"0818", X"0914", X"07B2", X"0567", X"026E", X"FE79", X"FE1A", X"FA03", X"F884", X"F995", X"FC33", X"FB8B", X"0164", X"0074", X"00CA", X"FCDE", X"FEE2", X"FEA3", X"FE2D", X"FFC4", X"0074", X"0392", X"01D1", X"026D", X"0444", X"0769", X"0611", X"0711", X"08A8", X"0525", X"FFF2", X"FDCE", X"FB33", X"FB62", X"FA40", X"F6C7", X"F7E1", X"F9E9", X"F96B", X"FC6E", X"FF03", X"023A", X"0154", X"FBE1", X"FC89", X"FDBC", X"FE3A", X"FF01", X"FFC6", X"02BC", X"0205", X"0365", X"05AC", X"05DE", X"04DB", X"04A0", X"02B3", X"FF5C", X"FC08", X"FAC5", X"FA4D", X"FABC", X"F952", X"F908", X"F95D", X"F936", X"F955", X"002A", X"0206", X"00AA", X"FDA2", X"FCCE", X"FF60", X"FF45", X"001C", X"02EB", X"0345", X"026A", X"0477", X"0535", X"030A", X"0070", X"0008", X"FE9D", X"FA04", X"FB27", X"FB58", X"FB28", X"FD22", X"FF79", X"FCA4", X"FB5E", X"FC19", X"F810", X"F5F6", X"FB00", X"FDCE", X"FF01", X"FBA5", X"FDDA", X"01B9", X"FEB5", X"01E2", X"03A7", X"0387", X"033A", X"00D3", X"0120", X"FF9B", X"FAF1", X"FA48", X"FACE", X"F9EB", X"FB82", X"FEC2", X"FF22", X"FF6D", X"FF30", X"FC86", X"FCE8", X"FE77", X"FA52", X"F530", X"FAC1", X"FE20", X"FF15", X"FFF3", X"FDC0", X"0035", X"01A2", X"000B", X"027B", X"FEC7", X"FEF4", X"FD76", X"FCAC", X"FBFC", X"F90E", X"FD06", X"FE5C", X"FCE0", X"FDCB", X"0235", X"0300", X"01EB", X"0254", X"FF72", X"0115", X"01EB", X"0103", X"FB12", X"FC2C", X"0059", X"0038", X"FB96", X"FE9B", X"FFB8", X"01C7", X"02DD", X"FEEA", X"FA87", X"FB59", X"FE96", X"FB9A", X"FB3E", X"FC66", X"FFDA", X"FFF5", X"FEA6", X"0179", X"023A", X"02C3", X"0243", X"0036", X"029E", X"0147", X"0552", X"053F", X"045B", X"0132", X"02EE", X"0077", X"FFD8", X"FE92", X"02B5", X"FEF0", X"FE05", X"FD8D", X"FD74", X"FCBC", X"FD35", X"FC83", X"FEFF", X"00F8", X"00DF", X"FF0D", X"FE56", X"0277", X"01A3", X"FFE7", X"FEFE", X"FCDA", X"0276", X"0418", X"092D", X"089E", X"0544", X"0688", X"043F", X"FE8A", X"FFD5", X"FE56", X"006F", X"FB04", X"FBB4", X"FE27", X"FC2E", X"FD39", X"FD92", X"000A", X"01F6", X"0077", X"FF48", X"FE38", X"FEF3", X"003A", X"FEDA", X"FF84", X"FC68", X"000B", X"019E", X"025D", X"0826", X"05F0", X"0585", X"082A", X"02C6", X"FF5B", X"FEE4", X"FBCD", X"FEAD", X"FD15", X"FCD1", X"FE21", X"FEF9", X"FCD2", X"FE5E", X"01DC", X"008F", X"FEC0", X"FD81", X"FDB9", X"FE30", X"0095", X"FECD", X"FF7E", X"0034", X"00C5", X"0100", X"016B", X"0439", X"07BD", X"0866", X"0326", X"01AE", X"005E", X"FFA5", X"00D9", X"01F6", X"0146", X"FDA4", X"FD4C", X"FC73", X"FC3B", X"FFB6", X"02C9", X"0226", X"FD56", X"FC92", X"FB30", X"FE56", X"FDF8", X"FDF0", X"FE8E", X"010A", X"006E", X"01BB", X"04DC", X"0620", X"08DF", X"0B0B", X"06B2", X"0325", X"0063", X"FF67", X"0027", X"03F1", X"0037", X"FCBC", X"FD88", X"FD7D", X"FDB5", X"FFE8", X"0268", X"00D8", X"FE9E", X"F94F", X"F8A8", X"FD9E", X"FE7B", X"FF03", X"00BA", X"0034", X"01D7", X"0257", X"0641", X"07AE", X"0999", X"09D4", X"0610", X"03C9", X"0236", X"FED8", X"FEE3", X"031D", X"01AA", X"012F", X"FE1A", X"00C2", X"004D", X"0263", X"0251", X"015D", X"FF2E", X"F8A7", X"FA35", X"FEFB", X"0030", X"0424", X"0367", X"04B6", X"0271", X"04BE", X"0774", X"07DF", X"0A9A", X"062E", X"014E", X"FE6B", X"FFB8", X"FF88", X"0021", X"0581", X"028B", X"02A9", X"02F0", X"03FB", X"0417", X"0414", X"03B2", X"0294", X"014F", X"011C", X"FFCC", X"FF11", X"00F8", X"0152", X"0299", X"033A", X"044F", X"0552", X"0A82", X"0843", X"0A32", X"04ED", X"0214", X"FD39", X"0012", X"012B", X"016D", X"04E7", X"07CE", X"0709", X"0573", X"029F", X"05AD", X"0574", X"0454", X"00AD", X"0233", X"028E", X"0027", X"00DE", X"004D", X"00B0", X"00E4", X"02DD", X"04F4", X"041D", X"061E", X"07B7", X"0830", X"077D", X"0087", X"FF19", X"FF3C", X"0015", X"0538", X"079A", X"0549", X"04EA", X"060E", X"04A5", X"044E", X"053C", X"0319", X"01AC", X"0342", X"03A7", X"02A0", X"0174", X"0188", X"FF95", X"00AC", X"01C2", X"01D5", X"0413", X"034C", X"04B2", X"0543", X"0247", X"0413", X"FEE0", X"0024", X"FFB7", X"02C0", X"04CD", X"04C3", X"041A", X"0492", X"040B", X"023C", X"00FA", X"0220", X"0097", X"01B0", X"01D7", X"0069", X"FFA6", X"0090", X"FEA5", X"FD19", X"FD74", X"FF68", X"0045", X"0197", X"03A1", X"01AD", X"0079", X"FDD7", X"00BB", X"FF70", X"0030", X"013D", X"05F7", X"00B2", X"0137", X"0245", X"01B6", X"0070", X"FCC8", X"FFCE", X"FE2F", X"FEB5", X"FF02", X"FE50", X"FEC3", X"FE15", X"FD2B", X"FCE7", X"FCEA", X"FD9E", X"FE48", X"0303", X"02D3", X"0375", X"FE68", X"FCA4", X"FFA6", X"0061", X"FEFE", X"FFF6", X"03A1", X"0352", X"00F5", X"0242", X"036A", X"038B", X"FF22", X"FFB7", X"00C8", X"0162", X"0187", X"0026", X"0114", X"0377", X"0252", X"00D1", X"FEEE", X"0168", X"FEFB", X"FF4B", X"00C1", X"03EF", X"FE81", X"0041", X"00E3", X"FFAD", X"FED3", X"0083", X"FB54", X"FE07", X"00E4", X"022D", X"00BA", X"0190", X"01D3", X"0386", X"03D9", X"043E", X"0226", X"020A", X"0462", X"05DF", X"05F9", X"0508", X"071E", X"0565", X"04E9", X"0160", X"0042", X"0140", X"0272", X"00D5", X"0058", X"FF82", X"FFE9", X"0038", X"FFAF", X"FEFD", X"FE99", X"FF47", X"0001", X"0328", X"021A", X"0469", X"0381", X"030F", X"06D6", X"0844", X"056F", X"06CE", X"0848", X"09A1", X"06BE", X"072D", X"0678", X"0424", X"00DF", X"0292", X"FF6E", X"FFA7", X"FF6C", X"0139", X"FF6F", X"00C2", X"00DC", X"FFA3", X"FE3D", X"FE12", X"FEDA", X"FDE1", X"FD81", X"FDC2", X"FD31", X"FB5A", X"F91E", X"008C", X"FD8B", X"FEE4", X"FEAD", X"001B", X"FF80", X"01E1", X"0195", X"00C3", X"FD20", X"FFF0", X"0037", X"0119", X"FFE2"),
--        (X"003E", X"FF6E", X"00B3", X"FF2F", X"FF86", X"0002", X"008D", X"0024", X"FFC1", X"FEDE", X"FE71", X"0057", X"FF9D", X"015C", X"FFAA", X"018C", X"FF8C", X"0082", X"01AE", X"FFB6", X"0037", X"0020", X"FEFE", X"0072", X"002E", X"00D4", X"FF97", X"012B", X"FFCB", X"FEED", X"00C3", X"00B4", X"FF56", X"FF6A", X"FF32", X"FD9F", X"FE45", X"FD89", X"FD50", X"FBCF", X"FBBE", X"FD3F", X"FFBB", X"0043", X"FFE5", X"FD4F", X"FD51", X"FD73", X"FCE1", X"FE3A", X"FF07", X"FF87", X"0037", X"004F", X"FFE3", X"FFF4", X"FF85", X"FFBE", X"FF13", X"FFB1", X"FEF3", X"FF06", X"FC59", X"FCF6", X"FCAE", X"FCD5", X"FC84", X"FBD3", X"FB4D", X"FA90", X"FA1F", X"FD42", X"FB88", X"F876", X"F871", X"FB7D", X"FC2D", X"FC94", X"FD5F", X"FF55", X"021B", X"0318", X"FEAE", X"003B", X"FFF5", X"FFAA", X"0194", X"FFE8", X"FE35", X"00DD", X"FF63", X"0189", X"FF6C", X"01A7", X"00B6", X"0248", X"011D", X"0005", X"FE56", X"FDE8", X"FAA2", X"F8C9", X"F86A", X"F713", X"F9C5", X"F9E6", X"FAA8", X"FDEC", X"009F", X"0393", X"FE96", X"012B", X"FF42", X"FEAC", X"040B", X"03AC", X"FF3B", X"0196", X"02F5", X"01CD", X"0492", X"06B3", X"059A", X"0335", X"04C3", X"02B4", X"00A7", X"FFB2", X"FF6B", X"FC79", X"FC0B", X"FB08", X"FB30", X"FAA2", X"FA14", X"F87C", X"FC90", X"02F2", X"011D", X"FF8F", X"011B", X"007C", X"031A", X"0330", X"01D7", X"0392", X"FF12", X"0190", X"01CB", X"0262", X"009B", X"02BE", X"0323", X"038B", X"01AE", X"01F2", X"FF15", X"FF9D", X"FDED", X"FF2B", X"FE3A", X"FEAB", X"F9DF", X"F815", X"FB58", X"007D", X"0009", X"FF09", X"FECE", X"00E6", X"02AD", X"05DC", X"0279", X"FF8B", X"00C4", X"FE52", X"FE6E", X"0150", X"02DE", X"0587", X"049E", X"060F", X"05F7", X"0651", X"05C7", X"0518", X"0305", X"0398", X"02C8", X"0118", X"FAFC", X"F6C3", X"FA51", X"01D3", X"FF72", X"FE5E", X"FFFC", X"0271", X"0297", X"03D0", X"02B1", X"FE83", X"004A", X"FDFB", X"FF4B", X"012E", X"0308", X"05B1", X"05BE", X"0805", X"055F", X"059F", X"04EF", X"0335", X"03D2", X"03C5", X"04E9", X"0374", X"FFC8", X"F906", X"F8E1", X"FCDA", X"FFEF", X"FE0B", X"FD53", X"0364", X"0076", X"0406", X"01A6", X"018B", X"02C7", X"01D9", X"011A", X"0156", X"03A3", X"03DD", X"04BC", X"0559", X"0677", X"0558", X"0218", X"03D3", X"0296", X"028A", X"016D", X"00CC", X"010C", X"FBD6", X"FBF5", X"FD8E", X"015A", X"0109", X"0099", X"027D", X"FF67", X"0513", X"03C7", X"063C", X"05BA", X"02AC", X"016A", X"01FB", X"0342", X"0569", X"0343", X"05A2", X"0659", X"0541", X"0079", X"00CA", X"0038", X"FEAA", X"FECA", X"FF13", X"019A", X"FDE6", X"FD1A", X"FEC6", X"02D2", X"01EC", X"019B", X"02C9", X"0594", X"067C", X"02FA", X"034D", X"0642", X"01A8", X"0019", X"FFFC", X"00C5", X"0037", X"00E7", X"0369", X"07A1", X"0112", X"FEFE", X"FEF3", X"FEA2", X"FF38", X"0024", X"0024", X"FE8C", X"FF46", X"FD73", X"FEBE", X"033C", X"02AF", X"00EE", X"015B", X"05CB", X"054E", X"055F", X"0381", X"014B", X"FE88", X"FF1A", X"FD9D", X"FE32", X"FEDD", X"FDE0", X"025B", X"0751", X"020D", X"FE93", X"0102", X"023F", X"0171", X"0281", X"FFBC", X"FFE8", X"FFA0", X"004D", X"0225", X"0474", X"0253", X"00B1", X"0307", X"0668", X"0255", X"05CC", X"0213", X"FCDF", X"FF3B", X"FD5B", X"FCDD", X"FB29", X"F84A", X"F8A8", X"FFF2", X"07C8", X"029C", X"0076", X"012B", X"0385", X"0391", X"00DC", X"0029", X"FD91", X"FCCB", X"FEA7", X"04C7", X"0964", X"05CA", X"FEB8", X"021F", X"0525", X"03B6", X"03D2", X"FCA6", X"FC4A", X"FD03", X"FC56", X"FB0A", X"FA13", X"F84A", X"F992", X"00DD", X"05D0", X"01A4", X"00DF", X"029D", X"00CC", X"FFFE", X"FF1B", X"FEEF", X"FD3B", X"FCE7", X"FF13", X"0471", X"09D5", X"0370", X"FE9A", X"0031", X"015C", X"030E", X"00AF", X"F9A7", X"FB90", X"FCA1", X"FB44", X"FBE1", X"F7E6", X"F80F", X"FAB8", X"026E", X"0486", X"019E", X"FF1A", X"0188", X"FF87", X"FF82", X"006C", X"FD75", X"FF72", X"FEDB", X"FD3A", X"02D4", X"0AE4", X"0271", X"FF67", X"0154", X"FE8D", X"0088", X"FE6F", X"F9C3", X"FD61", X"FCD7", X"FD48", X"FC05", X"FC39", X"F924", X"FE8C", X"02A1", X"00C1", X"FFBC", X"FFCA", X"FF01", X"0214", X"FFF4", X"FF90", X"0116", X"0075", X"FEB6", X"0064", X"0411", X"0999", X"02B5", X"011C", X"0045", X"042A", X"01F9", X"00C5", X"FC44", X"FCF2", X"FFAF", X"FD2E", X"FE1D", X"FDED", X"FD62", X"00E4", X"00A1", X"FF52", X"FDA1", X"0073", X"021A", X"000B", X"000F", X"FEBC", X"018F", X"027B", X"0157", X"0095", X"049B", X"0A7B", X"039C", X"008D", X"0281", X"006B", X"041A", X"016D", X"FD26", X"FC30", X"FD22", X"FDCB", X"FF47", X"FE08", X"FE97", X"01E7", X"0058", X"FD30", X"FF16", X"FF75", X"FF82", X"FD98", X"FFE3", X"FFC2", X"0104", X"02FB", X"01D1", X"0295", X"0500", X"077E", X"025C", X"0273", X"002F", X"015D", X"036B", X"00D4", X"FE38", X"FDED", X"FDB5", X"FE31", X"FED1", X"FF1A", X"FC50", X"FCA1", X"FDE0", X"FF16", X"FEB9", X"FEC1", X"FEC4", X"FFA6", X"FFB3", X"FF02", X"00D1", X"034C", X"03AA", X"0130", X"059D", X"06C6", X"0128", X"FEC7", X"FEFB", X"00B5", X"009D", X"0107", X"FF8E", X"000A", X"00EE", X"FFA1", X"FDDA", X"FC98", X"FCC7", X"FCBF", X"FE47", X"FDC2", X"FD52", X"FE2E", X"FE21", X"FFA8", X"007B", X"FFA8", X"0194", X"02F4", X"0310", X"0302", X"07AF", X"0536", X"02B5", X"FF7D", X"FD5D", X"FFDD", X"0032", X"01A4", X"027C", X"02C8", X"0144", X"0174", X"FE4D", X"FB46", X"FA43", X"FB8A", X"FD8B", X"FC69", X"FC87", X"FEC4", X"FEF2", X"FF85", X"0174", X"02A4", X"0234", X"0201", X"0562", X"04C3", X"0804", X"0308", X"000B", X"012D", X"00AD", X"01F1", X"010C", X"0159", X"049C", X"0579", X"0445", X"02E3", X"0004", X"FCD0", X"FC07", X"FC7A", X"FE55", X"FF25", X"FD23", X"FDF7", X"FED2", X"FFE8", X"004A", X"00F8", X"FDD5", X"0059", X"0228", X"057F", X"037D", X"FDB5", X"FF47", X"FEF2", X"008F", X"030D", X"01A6", X"038D", X"0541", X"074B", X"0659", X"0329", X"03E2", X"00E9", X"FEBD", X"FF72", X"FCD9", X"FF08", X"FEE2", X"FDEC", X"FDE6", X"FD0F", X"FD53", X"FEE2", X"FDAA", X"FF2A", X"023C", X"05DE", X"0364", X"FBFA", X"FEA9", X"FFE3", X"FF73", X"0117", X"0357", X"0409", X"0517", X"03BD", X"02D7", X"0685", X"021E", X"023C", X"00EE", X"006F", X"FF3A", X"FDE2", X"FCF4", X"FD7D", X"FF07", X"FE56", X"FE99", X"000F", X"FF05", X"009A", X"0157", X"02E1", X"FF1C", X"FDF8", X"FEF2", X"FFAA", X"003A", X"01D8", X"016A", X"02EB", X"02C3", X"05E3", X"061A", X"06EC", X"0463", X"0446", X"0342", X"02B9", X"00E8", X"0023", X"0107", X"FFBB", X"00C4", X"00B1", X"0230", X"010C", X"02F8", X"00C6", X"0119", X"0127", X"FE1E", X"00D2", X"FF87", X"0184", X"011C", X"00B8", X"019D", X"0336", X"07DE", X"06F1", X"087B", X"0A1C", X"08B5", X"05EE", X"07C7", X"0880", X"0868", X"07B3", X"04C1", X"065E", X"0630", X"057B", X"04FE", X"06D3", X"0439", X"020A", X"009D", X"01F4", X"0122", X"00A4", X"FFE1", X"0009", X"FFDF", X"005E", X"0121", X"027D", X"0501", X"063C", X"09C6", X"0A9E", X"0B9E", X"0A0F", X"091A", X"0A29", X"0B4F", X"0E0B", X"09FA", X"0A10", X"0A73", X"0BF6", X"0930", X"070E", X"04B3", X"03A2", X"02B3", X"01F0", X"02AF", X"0068", X"0080", X"FF05", X"FF39", X"FF8E", X"FFA1", X"0068", X"00BD", X"0404", X"038B", X"041A", X"033B", X"050E", X"020D", X"0411", X"060F", X"08EC", X"072C", X"06D2", X"07FA", X"068C", X"04F3", X"027C", X"05DB", X"0498", X"02E4", X"0051", X"0064", X"FFD1", X"FF68"),
--        (X"0067", X"FEB0", X"0021", X"008D", X"00DA", X"FF78", X"0029", X"0095", X"FFE3", X"FF68", X"0095", X"FEC0", X"0069", X"006B", X"0181", X"FEF7", X"FEFA", X"0002", X"FEF5", X"FFFE", X"005B", X"FFC8", X"0005", X"0002", X"0082", X"0004", X"0181", X"FFC4", X"FE34", X"00AB", X"FF40", X"FFB5", X"00FB", X"0029", X"FF7A", X"FE23", X"FF32", X"FF03", X"FE6A", X"FCED", X"FDB5", X"FDC2", X"0278", X"0090", X"FCCB", X"FCAD", X"FEE5", X"0012", X"FFB2", X"00A9", X"012A", X"0075", X"FFC1", X"0006", X"007E", X"FF89", X"007D", X"FE61", X"FEE3", X"FEE6", X"FEDC", X"00AE", X"FE6E", X"FCA2", X"FC61", X"FDB2", X"FB89", X"FB47", X"FF2D", X"019D", X"0101", X"021C", X"0416", X"00A4", X"013F", X"00D1", X"001C", X"FF11", X"0020", X"FED2", X"FCEA", X"FDB2", X"FFCA", X"0012", X"0000", X"0082", X"01FC", X"00F0", X"0087", X"FC6D", X"FE23", X"FB88", X"FB7A", X"FF09", X"FFA1", X"FB2F", X"FD41", X"FDCE", X"FE55", X"0066", X"0120", X"0109", X"043C", X"0138", X"020B", X"0262", X"01FF", X"01F7", X"002D", X"0302", X"FEBB", X"00DD", X"0075", X"00ED", X"021F", X"00FB", X"FE7F", X"FBE2", X"F9E9", X"F8C7", X"F7E9", X"FA61", X"FBC6", X"FBCA", X"FCFA", X"FFC1", X"016E", X"03E6", X"005E", X"00EB", X"02BB", X"FFD5", X"0000", X"00C8", X"01AF", X"027D", X"01CF", X"0275", X"01C4", X"FE96", X"00B4", X"FF70", X"01CC", X"FFB6", X"FC17", X"FE6E", X"FABD", X"FACB", X"F4BB", X"F717", X"F769", X"FAA6", X"FA93", X"FD67", X"FAC4", X"FB69", X"FCC7", X"FDB7", X"FFF8", X"FFFF", X"0466", X"00FE", X"012F", X"FF0F", X"FF5D", X"0086", X"00F1", X"FE5F", X"0007", X"FF60", X"FE8F", X"00AD", X"003A", X"FD59", X"FCD7", X"F914", X"F6C2", X"F86A", X"F99B", X"FC68", X"FF21", X"0041", X"0152", X"0189", X"FF82", X"0160", X"03B0", X"03C3", X"03C1", X"01F0", X"FEC7", X"FE4C", X"0043", X"001E", X"00BB", X"018A", X"001C", X"FC69", X"FEAA", X"01B8", X"FE02", X"FD31", X"FD5E", X"FCF0", X"FA9E", X"F9E8", X"0023", X"00B7", X"0373", X"037C", X"043C", X"023B", X"0411", X"015B", X"0057", X"0159", X"0329", X"01F5", X"FEE1", X"00C0", X"FF2D", X"0316", X"FDFC", X"0001", X"FD60", X"00F2", X"FE7E", X"0037", X"FF2F", X"FE5B", X"FF0D", X"FD8C", X"FD59", X"FEA9", X"0017", X"0485", X"045E", X"03C8", X"02EB", X"0116", X"00ED", X"02DE", X"01E6", X"02B7", X"028E", X"0328", X"0110", X"01AE", X"0415", X"06F6", X"034B", X"03A2", X"FF22", X"023B", X"FEF7", X"0125", X"FE7E", X"FEF6", X"FEE9", X"FBCA", X"FE44", X"0053", X"03EC", X"0547", X"039F", X"0486", X"0380", X"0116", X"FE7D", X"01CB", X"0143", X"0149", X"FFA6", X"00AD", X"00A1", X"012E", X"0711", X"0B12", X"0830", X"03A2", X"FFC4", X"0347", X"0194", X"007D", X"008B", X"FF60", X"0070", X"FE2C", X"FF55", X"00D5", X"03F7", X"0588", X"0583", X"0551", X"0629", X"01F1", X"0046", X"0115", X"00A9", X"000E", X"FFA3", X"0217", X"008F", X"0516", X"0959", X"0C02", X"0771", X"0252", X"00C8", X"011A", X"060C", X"0248", X"0572", X"0269", X"FF25", X"0125", X"0127", X"0238", X"0391", X"03C3", X"0370", X"06ED", X"0719", X"05A3", X"02DA", X"01E8", X"040C", X"FFD1", X"0247", X"01B0", X"01DB", X"04C1", X"07AB", X"0AEF", X"088D", X"0276", X"003B", X"0262", X"0392", X"0617", X"0705", X"04AC", X"00E8", X"FFB7", X"FE0E", X"FDF1", X"FD58", X"FDB2", X"FD54", X"0324", X"055F", X"0318", X"02DE", X"0166", X"02AD", X"00F5", X"FF7A", X"FEE7", X"FCA0", X"FE4E", X"FD82", X"036A", X"064B", X"0314", X"00BE", X"0029", X"02B2", X"0712", X"0824", X"0205", X"FDF1", X"FBFD", X"FB58", X"FC95", X"F9F9", X"F785", X"F958", X"0176", X"0394", X"02B8", X"0167", X"FF91", X"FFFD", X"FFA2", X"FF6E", X"FB9D", X"F9B5", X"F7D6", X"F919", X"FF20", X"FD10", X"FD1E", X"01FA", X"0259", X"028F", X"0407", X"0446", X"FD47", X"FCBD", X"FA33", X"FC58", X"FA53", X"FA0D", X"F793", X"F9BB", X"FF38", X"0380", X"034F", X"FE91", X"FEEB", X"FEE6", X"FEDF", X"FE42", X"FB86", X"F9A3", X"F77E", X"F7D9", X"FA00", X"FB92", X"FE05", X"0269", X"0372", X"FD8D", X"0150", X"FEEB", X"FF4B", X"FF94", X"FC90", X"FD0F", X"FB84", X"FC65", X"FA0E", X"FA0C", X"015E", X"018F", X"00CF", X"FD66", X"FE62", X"00E0", X"FE87", X"FE0B", X"FBA4", X"F893", X"F783", X"F846", X"F88B", X"FC48", X"FD5C", X"0095", X"0149", X"FCBE", X"FFDB", X"0074", X"0148", X"017A", X"00C7", X"FE9D", X"FE70", X"FD53", X"FEF5", X"FB83", X"0023", X"FE06", X"FECA", X"FCD3", X"FC74", X"FF59", X"FD0E", X"FC38", X"F97E", X"F5BF", X"F4C6", X"F490", X"F35E", X"FBB8", X"FF3D", X"FF13", X"00ED", X"FAB7", X"FF7D", X"0009", X"FF66", X"026F", X"0138", X"FFF4", X"FFEC", X"FF56", X"FEDA", X"FEB3", X"FEB8", X"FF55", X"FF59", X"FCE1", X"FFE2", X"FEF0", X"FE46", X"FCFB", X"F8B2", X"F55B", X"F347", X"F554", X"F5AB", X"FD5B", X"FE07", X"0053", X"0004", X"FFD2", X"FD76", X"FF67", X"FEBB", X"00F5", X"FF04", X"FFEC", X"FFDE", X"FEE5", X"FFCB", X"FE81", X"012C", X"0125", X"FFB2", X"FDAF", X"0177", X"0189", X"0182", X"FD0C", X"F8E2", X"F373", X"F289", X"F3BE", X"FA4D", X"0068", X"FF3D", X"017A", X"003F", X"0388", X"FC68", X"FCF7", X"FE2C", X"FF80", X"FE8C", X"FF47", X"FF1D", X"FEB6", X"FCA6", X"FF6A", X"00A5", X"FE87", X"FD50", X"FEF2", X"00F1", X"0340", X"042D", X"FE44", X"F695", X"F3EB", X"F4B2", X"F7F2", X"FB6C", X"009E", X"0257", X"000B", X"FCAA", X"FE1D", X"FA63", X"FB17", X"FEA6", X"FEF7", X"FEF6", X"FEFD", X"FF71", X"FD30", X"FCA3", X"FC8B", X"FE94", X"FCE4", X"FBE3", X"001E", X"02B8", X"0130", X"00B0", X"FA5B", X"F5AB", X"F4BB", X"F5C6", X"F9F6", X"FE63", X"0089", X"00FC", X"FF47", X"FE9C", X"FB0D", X"F951", X"FBDA", X"FEDB", X"FF2F", X"01B9", X"0039", X"00A8", X"FE7A", X"FDDD", X"FFE6", X"FC86", X"FDEC", X"FDBF", X"FE72", X"FD78", X"FF49", X"FDB0", X"FAA5", X"F81D", X"F5CD", X"F52F", X"FA0F", X"FBED", X"FC3C", X"FF6D", X"FF41", X"FDF7", X"F9CB", X"F812", X"FCE1", X"FF18", X"0007", X"FE8B", X"FE47", X"FF52", X"FF14", X"0012", X"FE86", X"FE7B", X"004D", X"FF2D", X"FE4C", X"FD2D", X"FD19", X"F99C", X"FAA3", X"FA8C", X"F7D1", X"F94D", X"FC7C", X"FD05", X"FC08", X"0066", X"FF05", X"002B", X"FA10", X"FC01", X"FF59", X"0104", X"FEDC", X"FD96", X"FDD4", X"FD4C", X"FF35", X"FEAD", X"FF06", X"0003", X"FE59", X"FF23", X"FF81", X"FDBA", X"FBEB", X"F9B5", X"FB90", X"FEC4", X"FDD0", X"FDE9", X"FD26", X"FD76", X"FE47", X"FF43", X"0073", X"015B", X"FFFA", X"FE12", X"0125", X"0408", X"0397", X"00E6", X"0062", X"0109", X"0010", X"01A9", X"02B6", X"02CD", X"01A5", X"0110", X"007D", X"0087", X"001F", X"FF20", X"FF88", X"025A", X"FF58", X"FF63", X"FC0E", X"FCEB", X"FF24", X"001A", X"015A", X"FF38", X"FCFD", X"034C", X"04F2", X"076A", X"0591", X"06C9", X"097B", X"099E", X"0A90", X"0AA8", X"095E", X"05C8", X"075F", X"04DC", X"0617", X"05F6", X"071D", X"0813", X"0975", X"0AE9", X"06BD", X"01BC", X"0120", X"FE9A", X"FD8D", X"FF97", X"00BE", X"0117", X"0013", X"00A4", X"0244", X"0356", X"04EE", X"05D5", X"07FB", X"0ABD", X"0909", X"08B1", X"0833", X"09FA", X"0B4C", X"08A0", X"08EF", X"082A", X"0924", X"08C0", X"0A7E", X"0909", X"0741", X"016F", X"FECC", X"005A", X"FFF4", X"FEF0", X"011D", X"010D", X"000E", X"FFBF", X"00FB", X"00A4", X"02FD", X"0257", X"02B1", X"02CF", X"047C", X"047C", X"0391", X"0389", X"05F3", X"04D1", X"045E", X"0473", X"04C1", X"03FE", X"0345", X"02F5", X"04BC", X"0266", X"FF79", X"0135", X"006E", X"0077"),
--        (X"FFA7", X"0051", X"00AF", X"0188", X"FEA8", X"003F", X"0093", X"FF9A", X"FE00", X"0040", X"FFAB", X"0026", X"FE2C", X"FF55", X"FFEF", X"FECE", X"FEFD", X"006D", X"00AC", X"FFED", X"FE68", X"0015", X"FFAE", X"FF62", X"FF10", X"0195", X"FF14", X"FF6D", X"0059", X"0070", X"0005", X"FF89", X"FFEA", X"008F", X"FB77", X"FB2F", X"FC52", X"FB89", X"FCEE", X"FB55", X"FA17", X"F987", X"FF23", X"FACC", X"FB2B", X"FA12", X"FA9B", X"FB76", X"FBF7", X"FD25", X"FD02", X"FDE9", X"005F", X"00C1", X"FF4B", X"00D8", X"0093", X"FF04", X"FFBE", X"FD62", X"FE14", X"FE80", X"FA68", X"F994", X"F861", X"F81A", X"F5FA", X"F4A0", X"F5DE", X"F81D", X"F96A", X"F92A", X"FB02", X"FBBE", X"FC93", X"FB96", X"FAAB", X"FB40", X"FB4E", X"FBF8", X"FD8E", X"FF3B", X"FF86", X"011D", X"FFBA", X"0074", X"003E", X"FB9F", X"FDF0", X"FC4D", X"F96B", X"F791", X"F765", X"F489", X"F59C", X"F62A", X"F57B", X"F4E7", X"F69B", X"F90C", X"FA5C", X"FB4E", X"0022", X"FFEA", X"FED1", X"FFE4", X"FF93", X"FDBC", X"FE59", X"FEE1", X"FE14", X"003F", X"009F", X"FECE", X"0028", X"FDC8", X"00B3", X"FCB8", X"FB85", X"FCCB", X"FB9E", X"FB2B", X"FBD2", X"FF9B", X"0027", X"FE8A", X"FDC5", X"FE32", X"FFAF", X"006A", X"FE27", X"FD79", X"FE5C", X"00A0", X"FEAE", X"0170", X"060A", X"058F", X"0052", X"FD21", X"FFB4", X"FFB3", X"FDAC", X"FD63", X"FCC3", X"FD65", X"FE07", X"FF1B", X"FF4E", X"FDF1", X"FE00", X"01AA", X"0089", X"FEFD", X"FE06", X"FDE7", X"FD8A", X"0043", X"FC75", X"FE6F", X"FEE5", X"0050", X"FFA5", X"0027", X"0045", X"0109", X"FFA2", X"FF0C", X"FFF8", X"FF98", X"FE88", X"FBDE", X"FE2A", X"0034", X"00BA", X"015C", X"0165", X"016D", X"017E", X"FFE0", X"FDD3", X"FD77", X"FD91", X"FF1B", X"FE87", X"FF41", X"FF03", X"FE1D", X"0163", X"FDD1", X"016F", X"0024", X"0013", X"013F", X"0024", X"FFE0", X"FE4C", X"FEF5", X"0182", X"FF96", X"FC6E", X"0012", X"0011", X"01D7", X"04DD", X"0354", X"02D2", X"01ED", X"FF47", X"FBB4", X"FD41", X"FEAD", X"0141", X"02DA", X"0098", X"0091", X"FFC3", X"0051", X"0175", X"027B", X"060E", X"0436", X"FFEB", X"FF7D", X"FDAD", X"FE7E", X"FE61", X"FEE3", X"FC09", X"00D7", X"01C9", X"034B", X"0480", X"0367", X"0347", X"0378", X"0110", X"FE61", X"FB7E", X"FE2D", X"01CC", X"013A", X"025E", X"02A5", X"FFE7", X"017C", X"02F6", X"078C", X"0A16", X"0A90", X"052B", X"0430", X"017F", X"0070", X"FEC6", X"FBAD", X"FC92", X"0174", X"02D6", X"0257", X"03B3", X"0487", X"0558", X"062E", X"0646", X"FF2C", X"F8E0", X"FC84", X"FFF0", X"01FA", X"023B", X"0365", X"020F", X"0127", X"0237", X"053C", X"067C", X"0BD1", X"06AF", X"0078", X"0053", X"004B", X"00E8", X"FDFC", X"FFDE", X"FF26", X"03F9", X"0512", X"039C", X"0526", X"0606", X"06D3", X"07A1", X"02EA", X"FC80", X"FEFC", X"FF33", X"0046", X"002E", X"0137", X"FFB4", X"0035", X"016C", X"01FF", X"0479", X"06D9", X"05B5", X"02DD", X"FFD8", X"FEFF", X"0122", X"005D", X"0385", X"02C8", X"0419", X"0699", X"0738", X"0710", X"07C3", X"06FA", X"06FC", X"0436", X"FFA5", X"01D4", X"01CE", X"014D", X"FF91", X"FE7E", X"FE16", X"FC78", X"FC7C", X"FE21", X"0112", X"061F", X"06AC", X"0194", X"FD99", X"00AA", X"0184", X"02FF", X"0238", X"05DF", X"0706", X"0626", X"0397", X"04F0", X"063F", X"059E", X"0540", X"0316", X"FE24", X"FF7C", X"0360", X"007E", X"FEB0", X"FF04", X"FE95", X"003A", X"FE11", X"FCED", X"FD8A", X"01CB", X"0427", X"FF91", X"FFF0", X"01DA", X"00BC", X"02E1", X"0543", X"027F", X"03C4", X"0447", X"02E9", X"030F", X"016D", X"04E9", X"035E", X"FFD9", X"FEE8", X"0017", X"FFAC", X"00F2", X"0190", X"FFD2", X"0116", X"00CF", X"FE83", X"FB2C", X"FCA9", X"0254", X"0193", X"FD5D", X"0264", X"0015", X"01A3", X"FFBF", X"04C9", X"001E", X"0019", X"FFC8", X"FF1C", X"0004", X"0098", X"03DE", X"016B", X"FEFF", X"FF05", X"FF38", X"0180", X"03AD", X"0193", X"016B", X"0106", X"FD64", X"FD4B", X"FD38", X"FE22", X"0090", X"FBAF", X"FE37", X"0277", X"FFFF", X"FE2C", X"FF57", X"FF8C", X"FA29", X"FE43", X"FCF3", X"FF8C", X"016E", X"009C", X"01B8", X"01A8", X"FE4E", X"FE6E", X"FEE5", X"02B8", X"04EF", X"01CF", X"FF2B", X"FE7D", X"FE2B", X"001E", X"FF62", X"FDCF", X"FDDF", X"FE4A", X"FD3E", X"FFA8", X"FF54", X"FD92", X"FAD6", X"FC8B", X"FBB6", X"FEA2", X"FF7B", X"008D", X"0073", X"FFAF", X"0074", X"0268", X"FFB4", X"FFED", X"02EC", X"0421", X"03DD", X"FFF9", X"FDD7", X"FE3D", X"FEFA", X"FEF7", X"0146", X"FE8F", X"FB02", X"FCC9", X"FE02", X"006C", X"FE5D", X"FF82", X"FA50", X"FBB6", X"FDF6", X"FFD2", X"FF18", X"00F8", X"FFE4", X"FE61", X"0053", X"02BA", X"026E", X"00C1", X"0289", X"02A2", X"014D", X"FF37", X"FE88", X"FFFB", X"00D0", X"FDCC", X"01B6", X"0205", X"F759", X"FCDE", X"FBB3", X"002F", X"FF28", X"0016", X"FA70", X"FB2A", X"FDDF", X"FFD0", X"FF79", X"FE3E", X"FE50", X"FE0B", X"0053", X"FFBF", X"FEF6", X"FDC4", X"FDA8", X"FE6F", X"FC25", X"FBD8", X"0077", X"0219", X"FF62", X"FE37", X"00A3", X"FE4C", X"F6EF", X"FF4F", X"FCAD", X"FFD4", X"FFB6", X"FF12", X"FC4B", X"FCC6", X"FE90", X"0031", X"FD05", X"FAE3", X"FC44", X"FBA7", X"FC5B", X"FDD4", X"FBBF", X"FCA0", X"FCA7", X"FA5A", X"FB44", X"FD72", X"FD8E", X"0062", X"0057", X"FF37", X"FFE8", X"FF01", X"F826", X"FC63", X"FF63", X"002A", X"FEA5", X"FF17", X"F9D8", X"F97C", X"FCB8", X"FDDC", X"FC23", X"FB63", X"F9F6", X"FB4A", X"FB70", X"FC89", X"FCC9", X"F98C", X"FA07", X"FB94", X"FACE", X"FB5D", X"FEF7", X"FF86", X"00CA", X"01E8", X"030A", X"FF0F", X"FB62", X"FC18", X"012E", X"0051", X"FFB1", X"FC84", X"F907", X"FA10", X"FAB7", X"FCF8", X"FB44", X"FB72", X"FAC7", X"F97E", X"FBAD", X"FC43", X"FCC6", X"FC53", X"FA95", X"FCF8", X"FCBC", X"FA02", X"FBBA", X"01D2", X"024D", X"0263", X"01D1", X"FE55", X"FCC5", X"FB76", X"003C", X"FE8C", X"FEB7", X"FD62", X"FB35", X"FA90", X"F97D", X"FB40", X"FCE6", X"FC5B", X"FB1F", X"FB70", X"FEFC", X"01C2", X"017A", X"0067", X"FDD5", X"FD0C", X"FEE9", X"FDDC", X"FD14", X"FF0A", X"0249", X"01A2", X"0121", X"00A6", X"FFD2", X"0072", X"FFF3", X"0067", X"0053", X"FC05", X"FC99", X"F9FE", X"F935", X"FA4E", X"FB51", X"FE09", X"FC16", X"FED2", X"001C", X"0218", X"02BB", X"0153", X"030A", X"010C", X"FF15", X"000C", X"008F", X"FF2C", X"0131", X"FFDC", X"FF1A", X"FF4E", X"0217", X"FFA8", X"0079", X"FF55", X"0013", X"FCEF", X"FBDF", X"FB06", X"FC9D", X"FD3B", X"FF2A", X"027A", X"0227", X"038A", X"0282", X"0270", X"01BD", X"015C", X"01CD", X"0188", X"FE42", X"FEAA", X"0252", X"012C", X"FE31", X"FF80", X"FED4", X"FCD6", X"FC04", X"FD9E", X"FF98", X"FECC", X"FFA1", X"FF49", X"0196", X"022A", X"02EC", X"03B4", X"0769", X"093D", X"09E4", X"0AF5", X"0A8E", X"0666", X"05C2", X"075A", X"08E3", X"05D0", X"01A8", X"015F", X"FEBD", X"00FA", X"FFCD", X"0131", X"0356", X"01D8", X"FE58", X"FEDD", X"FFCE", X"FE99", X"FF21", X"FFB0", X"027E", X"03F1", X"0418", X"0605", X"059C", X"0571", X"0385", X"04D2", X"06D7", X"04C3", X"0449", X"05D6", X"0539", X"0183", X"FF20", X"FF2E", X"FE92", X"FF1A", X"001A", X"FED9", X"027F", X"FF3E", X"FFBD", X"FF98", X"00E4", X"0034", X"FE6E", X"FEFD", X"012D", X"FFC3", X"0096", X"FE77", X"00B0", X"017B", X"FFE4", X"0233", X"00B3", X"0136", X"01DD", X"FE76", X"01DA", X"01FE", X"01CD", X"0029", X"FF8B", X"FF67", X"00B2", X"016B", X"0099", X"FF3A", X"00D7", X"007C", X"0050"),
--        (X"0079", X"FF62", X"FFFC", X"FF68", X"00C2", X"FE27", X"0207", X"0134", X"FF51", X"0058", X"0041", X"0087", X"025D", X"01F7", X"0126", X"009C", X"FF7E", X"FDFA", X"FFFF", X"01C2", X"FE4E", X"FFDB", X"01C2", X"FFEB", X"FEBB", X"FF66", X"0023", X"FF51", X"FE82", X"FFB1", X"0060", X"FFB8", X"FFBC", X"FED8", X"00EB", X"01A3", X"04E8", X"0288", X"0440", X"0281", X"0312", X"02EB", X"FFC2", X"04CA", X"04E4", X"0415", X"0769", X"0595", X"0624", X"0556", X"02AB", X"0334", X"FF6E", X"005E", X"FFC8", X"0072", X"0006", X"FF8D", X"005E", X"0192", X"017D", X"01AE", X"02B2", X"0485", X"0382", X"0799", X"082D", X"08AA", X"0877", X"0874", X"0755", X"0ADD", X"0B11", X"0891", X"0741", X"04C8", X"061D", X"0871", X"07C9", X"050D", X"017A", X"0132", X"015C", X"FF4E", X"0000", X"018E", X"FF71", X"024D", X"0080", X"02FD", X"0517", X"03BD", X"032F", X"0688", X"0821", X"09FF", X"0D0F", X"0C88", X"0D1F", X"0C78", X"0A38", X"083D", X"0567", X"0464", X"016F", X"FF87", X"FF31", X"FF26", X"FE85", X"FFAA", X"01A4", X"00F0", X"009D", X"FFBA", X"00F4", X"0296", X"01DB", X"04A9", X"03DA", X"0293", X"0437", X"07A0", X"091E", X"041A", X"0544", X"08A2", X"06EB", X"0496", X"03A9", X"FF3B", X"FF8D", X"FE55", X"FC66", X"F9A0", X"F951", X"F89D", X"FA50", X"FCD9", X"0226", X"01B5", X"FF60", X"FF68", X"0171", X"0209", X"0445", X"0958", X"0805", X"0720", X"061F", X"0465", X"02F9", X"023F", X"030C", X"0105", X"FFA4", X"00EE", X"FF8D", X"FD2B", X"FD9E", X"FB8C", X"FB16", X"FB27", X"F8FB", X"F7D4", X"FB1E", X"FB16", X"00CE", X"010E", X"FFAD", X"02A8", X"00B2", X"058E", X"06C8", X"071D", X"0696", X"0533", X"049B", X"05E5", X"0127", X"010F", X"FEC0", X"FE3B", X"FE8E", X"FE64", X"FD72", X"FD57", X"FDCB", X"FD73", X"FE9A", X"FCC0", X"F8A8", X"F846", X"FA30", X"FAEB", X"FF1E", X"0151", X"FE93", X"0504", X"0387", X"07DC", X"09FE", X"05C1", X"04A8", X"02FB", X"0051", X"FFF4", X"FFF3", X"FF83", X"FEF5", X"FDD6", X"FC3D", X"FC4C", X"FC88", X"FF11", X"FEC5", X"0064", X"012B", X"FE80", X"FB2E", X"F7E3", X"F767", X"F890", X"FF55", X"FF9A", X"FCD3", X"0582", X"0394", X"093A", X"0A4D", X"03CF", X"02F2", X"001C", X"0048", X"FEE4", X"007F", X"0086", X"0121", X"0178", X"FF89", X"FE60", X"FD75", X"FDAD", X"02D0", X"02A5", X"01B5", X"FF20", X"FC99", X"F633", X"F570", X"F88C", X"FF1A", X"0037", X"0100", X"02F3", X"0469", X"090A", X"08E9", X"032A", X"00C5", X"00C6", X"FFA3", X"001B", X"FCEB", X"FE33", X"FFED", X"027D", X"056D", X"00DC", X"FFFA", X"0018", X"0056", X"011E", X"0178", X"FDDB", X"FDC1", X"FB3D", X"F69F", X"F9D7", X"FEFD", X"0238", X"FFC9", X"03BA", X"0691", X"0861", X"053F", X"01EB", X"03D9", X"0042", X"FFCC", X"FD0E", X"FDB5", X"FC90", X"FCFE", X"03D2", X"0546", X"0254", X"016F", X"00D4", X"0080", X"005D", X"00BB", X"FFB1", X"FE96", X"FE06", X"FAB9", X"FA66", X"FD06", X"0015", X"FFD7", X"04EB", X"091D", X"094E", X"06E2", X"01B9", X"0026", X"FEE5", X"FCB9", X"FD31", X"FB32", X"FA42", X"FA4D", X"010B", X"0220", X"0244", X"FFF4", X"FEB3", X"001C", X"FFF9", X"00C9", X"FF1C", X"FF5A", X"032B", X"FFCE", X"FB4F", X"FAD2", X"00DB", X"0102", X"0536", X"07B2", X"0423", X"044A", X"FF2D", X"FDC9", X"FF12", X"FF61", X"FDFA", X"F991", X"F887", X"F8BB", X"FBBD", X"01E2", X"00E3", X"0049", X"FF79", X"0097", X"FF38", X"FDF5", X"FDD4", X"FF42", X"025B", X"0523", X"0408", X"0280", X"03F7", X"FF94", X"01AB", X"0571", X"0328", X"FCE8", X"FA2A", X"F9B9", X"FB0E", X"FB2D", X"FA53", X"F996", X"F7F0", X"F961", X"FD61", X"0261", X"0041", X"01C5", X"0166", X"01C5", X"FE93", X"FD44", X"FE2E", X"0070", X"0558", X"0790", X"082A", X"0758", X"0233", X"FEE4", X"01AF", X"06B8", X"FE8E", X"F935", X"F681", X"F448", X"F604", X"F915", X"F8F5", X"F91B", X"F9ED", X"FA99", X"00C9", X"02B5", X"0361", X"0206", X"0144", X"013D", X"01D7", X"FFB6", X"022A", X"03F6", X"0771", X"067D", X"05BA", X"0590", X"039D", X"FFC4", X"0169", X"0562", X"FFDA", X"F3FB", X"F859", X"FA70", X"F63B", X"F671", X"F753", X"F88F", X"FDCB", X"FD6D", X"04BC", X"0648", X"036E", X"0231", X"00F2", X"0287", X"02AB", X"02D5", X"04BB", X"04B5", X"02DC", X"0465", X"040B", X"FF73", X"0256", X"0273", X"02C9", X"05E2", X"FE72", X"F6BC", X"F92F", X"FBDF", X"F9D1", X"F9C9", X"FBE7", X"FB81", X"FFDE", X"0439", X"04DA", X"0447", X"0085", X"00CB", X"FFB0", X"005D", X"03DC", X"025C", X"048B", X"023A", X"FF66", X"01D2", X"0652", X"03A0", X"0166", X"FEEB", X"0309", X"089A", X"01EC", X"FA9B", X"FA98", X"FB06", X"FC3B", X"FC34", X"FB24", X"FF34", X"0408", X"03B4", X"0296", X"026C", X"FF6A", X"FE56", X"004F", X"018B", X"01E3", X"00F9", X"0224", X"0457", X"FFDE", X"0101", X"098D", X"0372", X"FFB6", X"0141", X"00B2", X"070F", X"03D5", X"FC5B", X"FB21", X"FC66", X"FBD6", X"FD3B", X"FC42", X"00BF", X"040E", X"0313", X"0143", X"002D", X"FFD7", X"00C8", X"02B8", X"FFFF", X"01EB", X"FF45", X"023A", X"0332", X"015E", X"FD79", X"0661", X"0535", X"0437", X"0012", X"009E", X"0128", X"0747", X"0100", X"FD07", X"FBEA", X"FDB1", X"FC86", X"004D", X"038E", X"0509", X"03F1", X"012E", X"0164", X"031D", X"020A", X"01EA", X"0126", X"0153", X"FF63", X"0087", X"006B", X"FE09", X"FE2E", X"0400", X"0564", X"0207", X"00DE", X"FF01", X"0215", X"0916", X"04BA", X"FDA1", X"FFE7", X"FF73", X"FEBC", X"0124", X"01D6", X"03A9", X"01EF", X"0165", X"01D9", X"0233", X"019B", X"02D2", X"0393", X"00EF", X"02EB", X"0001", X"FCAC", X"FCF3", X"FF8B", X"0055", X"0406", X"0063", X"FFC9", X"0132", X"0314", X"0740", X"04F0", X"03DB", X"0145", X"01BF", X"014A", X"FF3C", X"FF88", X"00E6", X"0025", X"00EB", X"0348", X"0243", X"02D5", X"02DB", X"02B3", X"0197", X"0000", X"FD18", X"FAE9", X"FCFB", X"FF60", X"0291", X"0238", X"FFD3", X"0073", X"0207", X"052A", X"0627", X"039E", X"06BF", X"04B7", X"03C0", X"017F", X"0304", X"FF97", X"FF07", X"FC54", X"FC7B", X"FDB9", X"0280", X"FFF1", X"0174", X"010A", X"01A2", X"FDD8", X"FB53", X"FA8C", X"F9C6", X"FC13", X"FE39", X"FD54", X"FFD5", X"000B", X"0089", X"02C2", X"0299", X"036A", X"0763", X"05CC", X"04C5", X"02D8", X"02FD", X"FF98", X"FF10", X"FF15", X"FF06", X"FD1A", X"FF9E", X"FEBC", X"0079", X"002D", X"0030", X"FBE1", X"F8CF", X"FAAE", X"FAD0", X"FC65", X"FE78", X"0012", X"0025", X"FF20", X"FF03", X"041E", X"027A", X"0316", X"03AB", X"0470", X"031C", X"0127", X"016C", X"0113", X"030E", X"0266", X"02EA", X"03BF", X"0151", X"FF7F", X"FF88", X"FD0B", X"FD27", X"F92C", X"F94E", X"FB4A", X"FA86", X"FFD8", X"013C", X"02D2", X"0199", X"010A", X"FF6F", X"FE9E", X"FEE3", X"0253", X"01E5", X"0350", X"02D5", X"0723", X"0480", X"0109", X"028B", X"0686", X"01EC", X"01DB", X"FEC0", X"FD4F", X"FD4C", X"FBAF", X"FB35", X"FA07", X"F749", X"FA2B", X"F9E9", X"FE31", X"FE82", X"018C", X"0111", X"0080", X"00C8", X"005C", X"FE4B", X"FCF9", X"FFB4", X"0039", X"01C3", X"01CA", X"0120", X"0181", X"01C3", X"FEEB", X"0091", X"FE98", X"00F0", X"017B", X"02CB", X"00E3", X"0269", X"FF34", X"FD3D", X"FD34", X"FEB9", X"FF95", X"00AD", X"FF11", X"00B0", X"FF2A", X"0029", X"FF92", X"0003", X"000B", X"019E", X"020C", X"0066", X"020E", X"02A1", X"0419", X"01C4", X"0199", X"06AB", X"03FB", X"03AB", X"069F", X"061E", X"0424", X"0426", X"FF0D", X"FE6D", X"FE0C", X"0035", X"FEE5", X"FEC2", X"FFE1", X"FF79"),
--        (X"00E9", X"FFCF", X"00BC", X"FFD2", X"FF4D", X"00EB", X"FFAD", X"0180", X"0015", X"FF54", X"0076", X"FFC5", X"0102", X"000C", X"0021", X"FFBE", X"001B", X"FFAD", X"FF79", X"FF36", X"FEF5", X"0067", X"00E9", X"0022", X"FFF9", X"0084", X"FFC1", X"FF85", X"FFEE", X"0030", X"FFB5", X"00EE", X"FEC9", X"0007", X"02DC", X"0327", X"00FF", X"011F", X"020D", X"00E1", X"03B4", X"034D", X"0166", X"041C", X"0616", X"0547", X"028B", X"02A6", X"0242", X"0437", X"0321", X"0340", X"FF1F", X"008D", X"001A", X"FF33", X"009E", X"000C", X"0008", X"01D1", X"0356", X"0100", X"015E", X"036B", X"032C", X"080D", X"08D7", X"07DE", X"06D6", X"05C9", X"08A3", X"084E", X"0791", X"076F", X"040E", X"0295", X"0420", X"07A6", X"0636", X"05C7", X"0417", X"02E0", X"0080", X"0031", X"FEB5", X"0086", X"FFE6", X"03C6", X"01A5", X"03E6", X"0417", X"0490", X"06C7", X"074B", X"0937", X"0A2A", X"0868", X"0A7D", X"0A18", X"077C", X"0808", X"0698", X"030E", X"0687", X"07A1", X"062A", X"0317", X"0355", X"02A1", X"FF8A", X"FED0", X"00DE", X"002D", X"006A", X"FE2B", X"02CF", X"01C2", X"0313", X"03C3", X"042B", X"055A", X"045E", X"0367", X"0176", X"0328", X"045C", X"021C", X"01C2", X"015D", X"0246", X"023D", X"0151", X"0067", X"FFEC", X"FEC3", X"FE7E", X"FC7A", X"FC00", X"FF74", X"0155", X"FF98", X"FF9F", X"0001", X"01E9", X"0278", X"0335", X"03D5", X"0408", X"0597", X"04AD", X"03F3", X"008A", X"00A6", X"006F", X"00F0", X"00EC", X"FFEE", X"00E0", X"0066", X"FDA7", X"FD6F", X"FF4B", X"FE27", X"FBC4", X"FC7A", X"FB49", X"FB09", X"0052", X"0083", X"01D9", X"001F", X"05A7", X"0562", X"0500", X"03EA", X"049D", X"031A", X"047D", X"035A", X"0282", X"0188", X"01C3", X"FFF3", X"0068", X"FF53", X"FEEE", X"0028", X"FDF6", X"FD9C", X"FE99", X"FF97", X"FA72", X"F750", X"F62E", X"F7C4", X"FAFD", X"FFF6", X"0177", X"01AB", X"05C5", X"050B", X"042C", X"0385", X"0257", X"013C", X"0252", X"0252", X"046C", X"031A", X"01B1", X"0137", X"FD9B", X"FE13", X"FEED", X"FDB5", X"FFBA", X"FF2E", X"FE26", X"FFA8", X"FE8F", X"FA47", X"F5EF", X"F984", X"FC45", X"0394", X"0330", X"0165", X"051B", X"066B", X"050D", X"00FB", X"01A2", X"0207", X"01D7", X"0391", X"050C", X"0548", X"0219", X"025F", X"00F9", X"000D", X"002A", X"0155", X"FFF5", X"FFE8", X"FEF1", X"FEF2", X"FDF6", X"F8DB", X"F704", X"F6A3", X"FC7F", X"FF67", X"0366", X"038D", X"0768", X"04E0", X"030D", X"018D", X"0022", X"FF60", X"00E4", X"023D", X"0289", X"0336", X"0477", X"059C", X"0595", X"035C", X"0346", X"0256", X"0184", X"007B", X"0021", X"FEC3", X"FD91", X"FA1F", X"F8FD", X"F7AB", X"FFDD", X"FF5C", X"03C6", X"05B0", X"0984", X"0380", X"0491", X"0077", X"FECB", X"FCBA", X"FD40", X"FDE8", X"FFEF", X"FF4B", X"043C", X"0654", X"0785", X"0797", X"0617", X"0352", X"0349", X"0385", X"01C2", X"004F", X"FD8F", X"FA77", X"F85E", X"F8A1", X"FE11", X"00B9", X"0665", X"0684", X"0AB0", X"0456", X"FE75", X"FABB", X"FAEB", X"FAE0", X"FAF3", X"FBF3", X"FD09", X"FB8A", X"FC90", X"FC4B", X"0145", X"0221", X"0291", X"02CE", X"00DD", X"0284", X"02EE", X"004C", X"FE94", X"FB34", X"F8EE", X"F78C", X"FE39", X"0236", X"03D3", X"05DE", X"076E", X"0107", X"FAA4", X"FA7D", X"F918", X"FA90", X"FAED", X"FD03", X"FC70", X"F86A", X"F785", X"F8FF", X"F9DC", X"FE9B", X"0074", X"0145", X"FE4D", X"FCEC", X"FD44", X"0009", X"FE5F", X"0323", X"014B", X"FD63", X"010C", X"FFA7", X"022C", X"061A", X"05A0", X"0040", X"FBD2", X"FC0F", X"FA50", X"F9C4", X"FB1B", X"FE6B", X"F8DE", X"F96A", X"F98B", X"F885", X"FAEB", X"FE07", X"FF4C", X"FFB6", X"FCE1", X"FBAB", X"FF0B", X"FF62", X"030F", X"082F", X"066F", X"0030", X"023D", X"FF8A", X"0163", X"040F", X"0438", X"01E2", X"FEB8", X"FE24", X"FE35", X"FC6F", X"FC6B", X"FC62", X"FC34", X"FB64", X"FB4B", X"FA33", X"FA93", X"FD55", X"FF54", X"0095", X"029D", X"0104", X"012E", X"0320", X"02F2", X"0518", X"054D", X"0531", X"013C", X"FED7", X"00ED", X"022B", X"0437", X"02A2", X"01B2", X"01A4", X"FF1B", X"FC18", X"FDB4", X"FC78", X"FD21", X"FCF5", X"FD9D", X"FC82", X"FBBA", X"FCAD", X"FEF4", X"03A6", X"020A", X"07F4", X"0666", X"039F", X"03A2", X"066A", X"0709", X"0740", X"030D", X"00CD", X"00B0", X"0174", X"03A0", X"0860", X"0518", X"03D2", X"021C", X"FE75", X"FD3E", X"FCEC", X"FC6E", X"FD1B", X"FC73", X"F9B3", X"FD10", X"FCCD", X"003B", X"016C", X"071B", X"06C8", X"0601", X"0384", X"01B9", X"040F", X"0A72", X"081B", X"0285", X"FF99", X"006E", X"0199", X"0758", X"0550", X"03F5", X"02F7", X"010D", X"FF33", X"FDE1", X"FCEE", X"FB45", X"FB23", X"FA77", X"FC99", X"FD61", X"FE81", X"033D", X"0382", X"05E3", X"055D", X"057C", X"0396", X"01DC", X"01D6", X"0B2A", X"0814", X"03D0", X"01CA", X"FF67", X"0489", X"08F9", X"070C", X"0251", X"00A6", X"0183", X"013C", X"0023", X"00AB", X"FEF9", X"FEF5", X"FE0F", X"FF98", X"015E", X"01F6", X"0496", X"02D0", X"02C3", X"0389", X"0384", X"044B", X"0092", X"007E", X"06C1", X"045A", X"0219", X"FF50", X"0311", X"0470", X"0BD0", X"056B", X"0065", X"016D", X"04CC", X"04A8", X"0415", X"05B5", X"0449", X"05BF", X"0472", X"0295", X"0211", X"0136", X"0109", X"026E", X"01EE", X"01D7", X"012C", X"FF1F", X"FDA7", X"0034", X"0330", X"0261", X"FF65", X"0026", X"02F5", X"025A", X"0AC5", X"0564", X"043B", X"02DC", X"0417", X"04A7", X"0598", X"04D8", X"04FB", X"03F5", X"03FE", X"0327", X"0182", X"FFAD", X"0033", X"00B0", X"007E", X"02F3", X"FE6F", X"FC71", X"FD5A", X"FF7E", X"012A", X"0105", X"FD4C", X"006A", X"017A", X"03E8", X"0710", X"043B", X"01B4", X"018D", X"023F", X"00CA", X"02C8", X"0329", X"00A0", X"0341", X"0443", X"00FD", X"009B", X"FFEA", X"FF34", X"0149", X"00FD", X"FF5A", X"FDAC", X"FB9D", X"000C", X"008C", X"042E", X"0536", X"0063", X"FE75", X"FFE3", X"03A7", X"0362", X"00BD", X"029C", X"01A1", X"FFBF", X"0146", X"FE77", X"FF9B", X"01D2", X"0048", X"FFBB", X"002F", X"0118", X"FFF3", X"FE35", X"FF41", X"003F", X"FFED", X"FDDB", X"FEFB", X"FE63", X"FFBE", X"FD77", X"FE02", X"FF98", X"FFF6", X"0052", X"0144", X"019B", X"02B0", X"02ED", X"030A", X"0270", X"FE0D", X"FEE9", X"FEC0", X"FF58", X"FF17", X"0072", X"FFCF", X"FE9E", X"FDC2", X"FEA3", X"FECA", X"00C6", X"FEDC", X"FDFD", X"FF4C", X"FAAE", X"FD81", X"FF6C", X"FBE3", X"FEFB", X"007B", X"0021", X"00FF", X"03DD", X"075F", X"04CE", X"05F3", X"039B", X"0161", X"0077", X"01C1", X"023D", X"01B0", X"0284", X"0335", X"0209", X"00ED", X"007C", X"FED8", X"FF1B", X"FE94", X"FD2D", X"FD6D", X"FC2E", X"FF11", X"011D", X"01B7", X"FFA2", X"00CB", X"0220", X"FEFE", X"FF56", X"0477", X"0675", X"05D3", X"0310", X"05B0", X"05D4", X"03D8", X"04EA", X"03E0", X"0328", X"02F0", X"0183", X"006E", X"FEE9", X"FED7", X"FFD9", X"FCB7", X"FD57", X"FE05", X"F906", X"FD74", X"FFC6", X"01FC", X"006D", X"FFD5", X"FFBD", X"0029", X"FED5", X"FE99", X"00D4", X"023A", X"02BE", X"0388", X"03DC", X"0195", X"005A", X"FF4B", X"0148", X"0214", X"02FA", X"0567", X"0329", X"04AF", X"04B1", X"FECA", X"0106", X"02D1", X"FF35", X"FFA5", X"0013", X"FF26", X"0047", X"FFC0", X"010C", X"0007", X"0125", X"FF75", X"0138", X"FFD4", X"0161", X"0260", X"0325", X"0263", X"0029", X"FFB0", X"068E", X"039F", X"004A", X"02DE", X"033A", X"00D7", X"02BA", X"023F", X"0319", X"02B2", X"0317", X"020F", X"00BC", X"FF99", X"FF51"),
--        (X"FEEF", X"009A", X"0018", X"00A3", X"0044", X"01CA", X"FF73", X"FFD8", X"01BA", X"007C", X"FEB4", X"FFCE", X"014C", X"FFF8", X"FFB8", X"0093", X"FF86", X"0058", X"0025", X"00C9", X"FF82", X"FFA4", X"FFAC", X"FF2F", X"011F", X"FF87", X"01DE", X"00C9", X"FF08", X"003D", X"0064", X"FFF3", X"FFBF", X"0068", X"0146", X"007B", X"0068", X"0022", X"013C", X"FEC1", X"FE2F", X"000D", X"0244", X"0305", X"0064", X"018C", X"0208", X"03C8", X"02CA", X"01FC", X"FFE4", X"0088", X"FF79", X"0003", X"00C8", X"FEDA", X"FF59", X"00D1", X"010D", X"FCF7", X"FE9B", X"FF5B", X"0215", X"00A3", X"0451", X"06AF", X"083D", X"05A2", X"04EF", X"06DE", X"0673", X"045A", X"0385", X"FFDC", X"FFAE", X"FF76", X"02A8", X"0268", X"0187", X"0333", X"02B9", X"016A", X"FF0B", X"FEF3", X"0019", X"FFC4", X"000D", X"FDCE", X"00CF", X"008B", X"0147", X"0324", X"0307", X"0632", X"02A9", X"01D4", X"FFCA", X"012A", X"FF74", X"FEF1", X"FDD2", X"FCF6", X"FD3F", X"FC88", X"FEB9", X"FFBB", X"FF97", X"FFFB", X"FFD3", X"FF15", X"FF07", X"FF5E", X"002E", X"00B3", X"0069", X"FEA3", X"017E", X"0204", X"FF74", X"00C6", X"0076", X"0057", X"FF79", X"FAE5", X"FE44", X"FEAA", X"FF0E", X"FEDB", X"FF5B", X"00C2", X"FE5E", X"FF81", X"0338", X"0181", X"FE4D", X"FE74", X"FC79", X"FB9C", X"0007", X"0371", X"001E", X"0134", X"01EA", X"FF20", X"01AE", X"FE15", X"FEEB", X"00ED", X"015B", X"FF5E", X"FFDD", X"FEE4", X"002A", X"FEFA", X"002F", X"FFA3", X"FEDE", X"FE3D", X"FE01", X"003B", X"FE9D", X"FE2A", X"FE10", X"FE7C", X"FEAA", X"FD2C", X"FDC7", X"02D9", X"FFBB", X"FF89", X"FE9E", X"00F1", X"FEB9", X"FE2C", X"FF21", X"02BA", X"00EB", X"00C5", X"FFE0", X"FF58", X"0061", X"FFDF", X"FE66", X"00D8", X"FF2E", X"FE8A", X"FD23", X"FE16", X"FD33", X"FE10", X"FE09", X"FCA9", X"F9D5", X"FC31", X"FC41", X"FE6B", X"0021", X"FD7A", X"03AE", X"003D", X"0237", X"FF79", X"FE63", X"039D", X"0205", X"00A1", X"FFDA", X"FFBF", X"FFDA", X"0060", X"FF5C", X"0266", X"008E", X"FEBF", X"FDEB", X"FEE8", X"FC38", X"FEE9", X"FEFD", X"FEA2", X"FC77", X"FA57", X"FE12", X"FD4C", X"FE9D", X"0009", X"030C", X"0456", X"02EF", X"0257", X"025B", X"0205", X"00BD", X"00F5", X"010C", X"009E", X"0000", X"0217", X"0200", X"01B8", X"0066", X"FE6E", X"FD8D", X"FC7A", X"FC0E", X"FCC7", X"FC40", X"FCF9", X"FB30", X"FB53", X"FD3A", X"FBD4", X"FFAA", X"01B5", X"018A", X"0487", X"03B7", X"02AD", X"01E7", X"015C", X"0050", X"008C", X"0261", X"0156", X"0260", X"0252", X"01E2", X"0305", X"01BC", X"011A", X"FDFF", X"FF3F", X"FE3A", X"FC8C", X"FA5F", X"FA7C", X"F4EE", X"F609", X"F980", X"FCBF", X"00AA", X"012C", X"00E2", X"032E", X"041E", X"048B", X"00CD", X"0178", X"FF65", X"02A1", X"0247", X"014F", X"0178", X"FE38", X"FEE8", X"FF4E", X"FFFC", X"0173", X"01BF", X"0092", X"FF97", X"FE42", X"FB06", X"F73E", X"F1C1", X"F163", X"F7C1", X"FE2F", X"018E", X"037B", X"04B3", X"03C4", X"023C", X"035B", X"0009", X"017E", X"015A", X"039F", X"01CD", X"FFB4", X"FD07", X"FCBF", X"FC51", X"FEAE", X"01DB", X"00ED", X"0267", X"02C5", X"037F", X"0439", X"01A7", X"FBA2", X"F647", X"F348", X"F77A", X"FF01", X"00B4", X"0391", X"05C3", X"051B", X"0305", X"02D5", X"FF98", X"0086", X"0210", X"00E7", X"FE04", X"FD0E", X"FB91", X"FC04", X"FB5A", X"0087", X"02AF", X"04A2", X"033E", X"057C", X"069D", X"08CD", X"07E3", X"06A6", X"048A", X"FEB8", X"FAE5", X"01DB", X"0005", X"01E6", X"047A", X"0305", X"0176", X"FFB1", X"005B", X"FF3D", X"FEA8", X"FDC7", X"FD38", X"FB5C", X"FA74", X"FBFA", X"FF56", X"0490", X"04D4", X"0417", X"02E1", X"04E1", X"065C", X"0526", X"04F3", X"0630", X"0752", X"067C", X"01F3", X"02DE", X"FD90", X"FE24", X"0203", X"0186", X"0013", X"FFB5", X"0107", X"FE04", X"FC5F", X"FB1E", X"FB5F", X"FC41", X"FD58", X"00FB", X"02DC", X"035F", X"036C", X"0499", X"0230", X"023E", X"00AD", X"FE92", X"FFA5", X"FED9", X"FF30", X"0732", X"0606", X"013E", X"FF74", X"FD77", X"FF46", X"00ED", X"FC24", X"FC53", X"FDB9", X"FB6C", X"FBAC", X"FD20", X"0003", X"02D8", X"01A6", X"02B8", X"0489", X"03C3", X"02B5", X"02AD", X"011C", X"0033", X"F935", X"FA50", X"FCB1", X"FCF1", X"FCDA", X"05D1", X"06FF", X"023E", X"0126", X"FD75", X"FCB7", X"FFFD", X"FBA2", X"F928", X"FAFA", X"FD3D", X"00ED", X"09E5", X"0AE4", X"0948", X"0655", X"0511", X"0597", X"0412", X"03CC", X"003B", X"FF6B", X"FC4E", X"FC56", X"F9FC", X"F8DD", X"FB2A", X"FCB8", X"0727", X"0647", X"0250", X"FFD0", X"FD46", X"FFFA", X"FCBF", X"F839", X"F498", X"F642", X"FAB7", X"04D6", X"0B4E", X"0EE3", X"0A62", X"089C", X"06EA", X"070F", X"03EE", X"0155", X"FE19", X"FE13", X"FD3A", X"FD05", X"FC16", X"FABB", X"F99D", X"FC2B", X"08AC", X"0759", X"FF9E", X"022E", X"0002", X"FEFB", X"FD9D", X"FA22", X"F59F", X"F531", X"F8D8", X"001D", X"0729", X"07BF", X"04C1", X"03C9", X"03E0", X"046A", X"0286", X"FF52", X"FF37", X"FF20", X"FEC3", X"FF81", X"FD4D", X"FB7F", X"FC2F", X"FFAD", X"0A84", X"05F0", X"0358", X"FFAC", X"FEC0", X"FE4D", X"FA76", X"FAD9", X"F86E", X"F88F", X"F932", X"FC43", X"00AE", X"012A", X"00BA", X"FF43", X"00B3", X"008A", X"FF91", X"014A", X"FFAF", X"FFE6", X"0005", X"FF05", X"FE3B", X"FD3E", X"FC18", X"0073", X"09E9", X"04B1", X"0356", X"00F6", X"FCB8", X"FD1F", X"FA9C", X"FB4B", X"F8C4", X"FA85", X"FB50", X"FBA8", X"FC6E", X"FF33", X"FF08", X"FF83", X"FF0D", X"FFF1", X"00FE", X"00C7", X"0084", X"0130", X"0162", X"0157", X"FE80", X"FC24", X"FDC6", X"03AD", X"079C", X"02E5", X"FFC1", X"00E9", X"0051", X"FB25", X"FBA6", X"FB4C", X"FCD3", X"FC88", X"FE0C", X"FDA5", X"FDAC", X"FEC5", X"FED4", X"FECA", X"FEDF", X"FFF9", X"FEE0", X"0147", X"0128", X"00AE", X"00EA", X"FEFD", X"FE45", X"FE24", X"FE9C", X"08E4", X"07D5", X"015C", X"0078", X"0078", X"00B7", X"FBEB", X"FCB8", X"FF3E", X"01C7", X"FFDA", X"FF77", X"FFEC", X"FD65", X"FE33", X"FE18", X"FE8B", X"FD59", X"FEBA", X"0012", X"0030", X"017F", X"014A", X"0040", X"FE21", X"FF09", X"FE58", X"FF4E", X"02E1", X"04BF", X"0024", X"002E", X"002D", X"FEDF", X"FD16", X"F867", X"FBDF", X"FF2D", X"FFAE", X"FE84", X"FE68", X"FCF2", X"FD6A", X"FCCB", X"FF46", X"0023", X"00F2", X"FF06", X"FFE4", X"00B8", X"0192", X"004B", X"0188", X"0098", X"FEEE", X"00DC", X"FF5D", X"01C2", X"FE41", X"FE47", X"FF82", X"00A3", X"FF8A", X"F99C", X"FB8F", X"FD91", X"FDF7", X"FFB2", X"FF86", X"FF48", X"FD91", X"FDEA", X"FED3", X"FC73", X"FE88", X"006C", X"005A", X"002A", X"0068", X"01B2", X"009A", X"00DD", X"FE0A", X"FDCF", X"FEB6", X"033F", X"01EE", X"0077", X"007D", X"FEF0", X"FDA4", X"FED6", X"FF8E", X"FDEA", X"FD59", X"FF42", X"FF5B", X"FECE", X"FF34", X"FE62", X"FEEF", X"FF7A", X"02F8", X"FF78", X"FEE9", X"FEE2", X"FF86", X"FFAC", X"FE80", X"FEB0", X"FC71", X"FC45", X"FAE2", X"FF69", X"FFCA", X"FFE7", X"FFBF", X"FF74", X"00BE", X"00C1", X"001A", X"FF40", X"01E6", X"0447", X"0730", X"0594", X"0226", X"00A3", X"00FA", X"003F", X"01D8", X"00E8", X"0108", X"FFAA", X"014A", X"FF5B", X"FCAB", X"FEBA", X"FECB", X"0120", X"FEF5", X"FF9C", X"00E2", X"005D", X"FF7A", X"002A", X"00B5", X"0067", X"005A", X"015D", X"FFE6", X"0209", X"0185", X"0189", X"FFB0", X"FF74", X"0015", X"02FD", X"039E", X"030C", X"0247", X"02AA", X"02D6", X"0407", X"026D", X"0396", X"02D4", X"018E", X"FF96", X"FFDA", X"FFA4", X"FFF6"),
--        (X"FFF2", X"0206", X"FF72", X"FFB5", X"FFBB", X"FF38", X"0222", X"0176", X"FFE4", X"FEF9", X"FFD8", X"0042", X"FFC1", X"00C0", X"0025", X"0034", X"FF3F", X"0034", X"011E", X"FE42", X"00D8", X"003D", X"000B", X"00E1", X"FFE8", X"FF77", X"0075", X"FF5A", X"01A0", X"FFB4", X"0185", X"0017", X"00A4", X"012B", X"0068", X"0155", X"0474", X"0326", X"0354", X"0307", X"052F", X"024C", X"00E0", X"013D", X"FD66", X"FE79", X"0566", X"0554", X"0574", X"0416", X"00BF", X"0072", X"FF11", X"0046", X"0011", X"FEE2", X"005E", X"0215", X"FF6B", X"FF0E", X"0086", X"024F", X"02AB", X"00A1", X"02EA", X"0206", X"04BB", X"04BB", X"0279", X"0113", X"FF4A", X"0229", X"02FA", X"02F5", X"0312", X"05BE", X"05C8", X"0524", X"07C8", X"04AD", X"02CF", X"FE6E", X"0105", X"000D", X"FFC7", X"00E4", X"FFF0", X"0115", X"02B4", X"0210", X"007D", X"0172", X"01EF", X"FE43", X"0071", X"FC7E", X"FCF6", X"FB45", X"FAB5", X"FEE1", X"FEE5", X"FE3B", X"04AA", X"010A", X"03F6", X"0535", X"078C", X"0B34", X"069A", X"FFA9", X"005A", X"0075", X"001E", X"FF98", X"FFE4", X"0194", X"0321", X"FF89", X"FE95", X"FED3", X"FF43", X"FC7E", X"FDD5", X"FDF2", X"FD0E", X"FD50", X"FF0F", X"FD6D", X"FDCC", X"FE7E", X"FFE4", X"01AB", X"0202", X"03C1", X"0209", X"07C6", X"052C", X"0393", X"05B8", X"037B", X"FFFE", X"002F", X"01D4", X"FF28", X"02F8", X"FE1E", X"FE52", X"FEFA", X"000D", X"FF9C", X"FEE9", X"FE5C", X"FF09", X"FF6E", X"FF9A", X"FD31", X"FD08", X"FD1A", X"FD13", X"00A8", X"0161", X"FE75", X"FFCF", X"02E4", X"0413", X"064C", X"06CC", X"03D5", X"FF2B", X"010E", X"FEE5", X"FE28", X"0085", X"FF57", X"FE5D", X"00D9", X"005E", X"0060", X"0076", X"01AC", X"02BF", X"FEE4", X"FF67", X"FF58", X"FDB1", X"FCFA", X"FB7B", X"FDA7", X"FF8F", X"FE01", X"FE7F", X"041A", X"0740", X"0B36", X"08CE", X"02DD", X"FFF7", X"FCED", X"FCA1", X"FB8A", X"00D7", X"FF4C", X"FE50", X"02CA", X"016B", X"FF8D", X"FF2E", X"FE22", X"FE5C", X"FE1F", X"FDE0", X"FF24", X"FDA5", X"FAD0", X"FD63", X"FB96", X"FD05", X"FEC9", X"FBD9", X"006B", X"05FB", X"08D0", X"09B7", X"03BB", X"FEA9", X"FBC8", X"FD37", X"FF59", X"FEE6", X"0069", X"017E", X"01A8", X"00BC", X"0120", X"FEC8", X"FEBC", X"FF6B", X"FF37", X"FBD3", X"FB63", X"F986", X"FA8A", X"FAD1", X"FAD1", X"FC38", X"FEA6", X"FD07", X"FD34", X"0739", X"0A31", X"0943", X"0208", X"FEC3", X"FC96", X"FE0D", X"FE26", X"0194", X"00E1", X"03EB", X"04DD", X"026C", X"0021", X"FF41", X"FE47", X"0030", X"0169", X"FDD0", X"F6FB", X"F5A9", X"F70A", X"F7A8", X"FA2E", X"FD1F", X"FE48", X"FEB1", X"01FB", X"03B9", X"0959", X"070C", X"0288", X"FF30", X"FE25", X"FD19", X"FEBE", X"02B7", X"0110", X"033F", X"043B", X"02E7", X"001F", X"01E9", X"0028", X"035D", X"0382", X"0359", X"FBE5", X"F55C", X"F65C", X"FA43", X"FBFC", X"FC70", X"FE55", X"FE4A", X"01E6", X"0489", X"069C", X"060B", X"023E", X"FFCB", X"FDBD", X"FDC7", X"FE20", X"00FE", X"0184", X"02F1", X"04AD", X"02CE", X"033B", X"0473", X"0460", X"0654", X"0B3F", X"0D35", X"04A6", X"FCFA", X"F9D8", X"FB05", X"FC7C", X"FDEA", X"FF45", X"00A9", X"046F", X"05F3", X"0703", X"0619", X"01FE", X"003A", X"FE2D", X"FA93", X"FDC1", X"019B", X"0464", X"05A3", X"05DE", X"0204", X"05CB", X"040A", X"0557", X"0686", X"0985", X"0BBC", X"07D1", X"006A", X"FD36", X"FE9E", X"005C", X"020A", X"02D4", X"0376", X"033B", X"0490", X"0275", X"02A2", X"FF73", X"FF98", X"FE51", X"FB36", X"FD6F", X"0030", X"0295", X"042C", X"030D", X"026D", X"0347", X"01B0", X"02D4", X"0438", X"081F", X"0866", X"0855", X"041E", X"00F2", X"0113", X"0262", X"03C1", X"0307", X"03BF", X"03DB", X"00C3", X"FF23", X"FC49", X"FD73", X"FFF1", X"006D", X"FD35", X"FAF8", X"FB63", X"FE3F", X"0145", X"0173", X"0470", X"0555", X"02D2", X"03F8", X"05A6", X"03D4", X"0469", X"066C", X"03D0", X"023A", X"0069", X"0082", X"002A", X"0197", X"0219", X"0054", X"022A", X"FD48", X"F8B4", X"FCF4", X"00E1", X"01F0", X"FF8F", X"F9F3", X"F744", X"F712", X"FAAA", X"0011", X"0271", X"04B3", X"0583", X"0611", X"058A", X"0558", X"0837", X"05DE", X"038F", X"014C", X"FEF1", X"FD1C", X"FD13", X"FEC9", X"0024", X"0206", X"FD59", X"FCCD", X"F70A", X"FACA", X"FFDF", X"0099", X"FF31", X"F8A7", X"F443", X"F5A1", X"F633", X"FC27", X"0142", X"0473", X"03B6", X"059D", X"063F", X"0622", X"093C", X"0409", X"015A", X"FE9B", X"FED2", X"FE3F", X"FC09", X"FE1E", X"02D8", X"0164", X"FE54", X"FB57", X"F79E", X"FD37", X"FE84", X"010B", X"FE68", X"F723", X"F36E", X"F5E1", X"F953", X"FB31", X"FD2E", X"FF64", X"0064", X"025C", X"0382", X"0500", X"04EB", X"0399", X"FF19", X"FEC2", X"FE1A", X"FEE9", X"FF79", X"010B", X"01E2", X"01A4", X"FE08", X"F834", X"FA9D", X"FB1B", X"FD22", X"0098", X"FF0D", X"F8A5", X"F877", X"F8FC", X"FC8C", X"FAD0", X"F9B2", X"FAD6", X"FC52", X"FD1A", X"FE2C", X"FE8C", X"0237", X"0127", X"00C7", X"FD25", X"FF4F", X"FDEE", X"0083", X"FFAF", X"0050", X"00C6", X"FE41", X"F8AA", X"F8E6", X"FACF", X"00F6", X"FEE8", X"0020", X"FBC0", X"FA51", X"FD2D", X"FC71", X"FA69", X"FBC2", X"FBA3", X"FA7A", X"FA7F", X"FB05", X"FCFD", X"FDD2", X"00D0", X"00EB", X"0105", X"FFB4", X"FF10", X"FE50", X"FFF5", X"0293", X"0160", X"FEB5", X"F8CE", X"FA5E", X"FD7F", X"FF22", X"FF37", X"FFBE", X"0036", X"FDF0", X"FCE0", X"FEBD", X"FD9A", X"FE1C", X"FBEE", X"FD5A", X"FB75", X"FB58", X"FF07", X"0150", X"018A", X"0278", X"0126", X"00AD", X"FEDE", X"FF5C", X"00FD", X"01F0", X"FF3F", X"FD21", X"FB00", X"FB5F", X"014B", X"0002", X"0059", X"03B4", X"02CD", X"008D", X"00B4", X"FF8D", X"FF5E", X"FF78", X"FEB9", X"FF38", X"FD88", X"FD66", X"FF2F", X"009E", X"0350", X"00DF", X"022E", X"FE68", X"FD4E", X"FED2", X"FE22", X"FE01", X"FD79", X"FB98", X"FB58", X"FE4C", X"0027", X"002C", X"0023", X"00D1", X"0292", X"0395", X"FFBD", X"FF82", X"0101", X"0070", X"0044", X"00F7", X"FF65", X"FF92", X"00E2", X"FFF2", X"0198", X"0185", X"01B0", X"FFE1", X"FCF7", X"FC46", X"FE5D", X"FBA9", X"FEFE", X"FCAA", X"0120", X"039B", X"008D", X"0041", X"0092", X"01A9", X"04B0", X"032F", X"016E", X"00F8", X"0295", X"0470", X"02C1", X"006F", X"FEF6", X"FFFE", X"000D", X"01BA", X"0091", X"0398", X"00A9", X"FD94", X"0068", X"0043", X"FD8A", X"FBF0", X"00BD", X"FF50", X"00AA", X"02A1", X"0117", X"FFEB", X"0117", X"0170", X"03BC", X"FFDD", X"FB8C", X"FEC4", X"0045", X"03FD", X"0311", X"0402", X"0354", X"014A", X"0132", X"0183", X"00A1", X"023B", X"0045", X"FF60", X"FFCE", X"FFC7", X"FEC0", X"FD8B", X"0040", X"FCA1", X"FBF1", X"FDDC", X"014E", X"FFA6", X"FF0D", X"02B5", X"FE45", X"FB43", X"FB94", X"FF08", X"00F1", X"FF15", X"00E8", X"020E", X"00DB", X"0069", X"FDF9", X"FF10", X"FDBD", X"FF17", X"014A", X"004F", X"01BB", X"028D", X"0040", X"021A", X"0515", X"031E", X"FDE9", X"FCBC", X"004F", X"FF58", X"FF69", X"0078", X"00F6", X"0253", X"FF54", X"FE9E", X"FD99", X"FDF1", X"FF75", X"FFDD", X"FD9C", X"0018", X"FEC5", X"FBF5", X"F822", X"FB21", X"FB02", X"FC0F", X"FB96", X"FDE0", X"FE99", X"FD80", X"0299", X"0111", X"010A", X"0056", X"0080", X"FFFA", X"00E6", X"FF6D", X"010A", X"FEF8", X"FDBA", X"FD8B", X"FF14", X"FDFC", X"FBB7", X"FDCD", X"0031", X"FF62", X"F968", X"FB2A", X"FB91", X"FBEE", X"FC59", X"FF85", X"FCFD", X"FD60", X"FC61", X"FAAF", X"FCE9", X"0226", X"00D1", X"FF7B", X"0123"),
--        (X"0090", X"FED6", X"00CC", X"FEBE", X"0041", X"0075", X"FFC4", X"FFE5", X"0097", X"FEB9", X"FEC5", X"FFAF", X"FFA3", X"0028", X"FF9A", X"FF97", X"007B", X"001F", X"002D", X"0101", X"0036", X"0162", X"FEA8", X"FF8D", X"FF17", X"0051", X"000E", X"FFBD", X"FF8C", X"FFC6", X"FEED", X"FFC6", X"0177", X"FF05", X"FBD9", X"FB24", X"FBF1", X"FC12", X"FD1E", X"FE77", X"FEBA", X"FD91", X"005E", X"FDB6", X"0087", X"FDA8", X"FDD5", X"F981", X"FB57", X"FDAE", X"FC6D", X"FF7E", X"0086", X"0093", X"01FC", X"0011", X"FF8B", X"FEEA", X"FF46", X"0165", X"00D5", X"FE2C", X"FBD7", X"F932", X"F5DC", X"F38A", X"F493", X"F67F", X"F786", X"F7A3", X"FA1F", X"F83F", X"FAAF", X"FD4C", X"FD44", X"FEB1", X"FE37", X"FCCF", X"FDD2", X"FBC2", X"FC09", X"FF79", X"FEE2", X"0132", X"FFC3", X"001B", X"FFDE", X"FC62", X"FF36", X"011E", X"FD43", X"FBC9", X"FBFE", X"FB23", X"FAA0", X"0051", X"FEB0", X"FDAB", X"00F5", X"FFB3", X"FFC7", X"FF9B", X"010A", X"FFF3", X"019B", X"010D", X"FE7A", X"FFCF", X"0217", X"FF00", X"0017", X"FF12", X"0036", X"001F", X"FFDB", X"0044", X"FEFA", X"FF2D", X"FFB2", X"00CE", X"FE6C", X"FFEB", X"000C", X"0200", X"01B0", X"0100", X"FFA7", X"FEC0", X"FFBA", X"0022", X"01BD", X"FFF2", X"FE50", X"FF42", X"FCBD", X"FBC5", X"01E0", X"04BC", X"0299", X"FFD3", X"FFD4", X"004D", X"FE50", X"0260", X"00A6", X"03AC", X"0333", X"02CA", X"043F", X"0162", X"0112", X"0356", X"0262", X"00F1", X"FEE4", X"FE37", X"FFAB", X"0058", X"FE7D", X"FE5F", X"FDB9", X"FB50", X"FC66", X"FB60", X"FAD0", X"00D6", X"0152", X"FE41", X"009B", X"FFE5", X"0176", X"02C1", X"FF9C", X"0680", X"059B", X"04FF", X"05BC", X"066B", X"0456", X"0311", X"024C", X"01C1", X"0015", X"0254", X"0319", X"040A", X"0178", X"00F9", X"FEDE", X"FECF", X"FE5E", X"0026", X"002D", X"01FC", X"0283", X"FED6", X"00B7", X"0020", X"0043", X"050F", X"04CF", X"06F0", X"06FC", X"0541", X"070B", X"0663", X"0261", X"013F", X"02F6", X"FFFE", X"00C6", X"0391", X"02C7", X"0351", X"034E", X"02F5", X"00CC", X"0242", X"0220", X"0329", X"05D0", X"047E", X"013C", X"0126", X"0040", X"FEF6", X"FFF3", X"06BF", X"03B3", X"0479", X"0550", X"0504", X"07AD", X"059E", X"027F", X"025A", X"0039", X"0198", X"012B", X"0237", X"0489", X"0378", X"05DF", X"0548", X"0324", X"03E8", X"0427", X"089B", X"0B48", X"08A3", X"04F9", X"03D1", X"003D", X"00A2", X"02C1", X"0228", X"04ED", X"044C", X"07DA", X"0533", X"05C0", X"03B2", X"0351", X"0155", X"0190", X"013B", X"FEE6", X"FF37", X"0182", X"0569", X"0646", X"0652", X"053A", X"0389", X"06E8", X"0B9C", X"0B68", X"07DD", X"04CB", X"FF3A", X"00F2", X"FFC7", X"0231", X"0721", X"04E7", X"03BB", X"0608", X"0418", X"041D", X"052D", X"0300", X"0270", X"0083", X"015A", X"FEE0", X"FF64", X"008C", X"01EF", X"0677", X"06DF", X"0532", X"0315", X"064A", X"0AEA", X"0B36", X"06C3", X"0656", X"0136", X"FEF2", X"FDF4", X"02CF", X"068C", X"0212", X"0395", X"0521", X"0355", X"0388", X"030C", X"049D", X"01F3", X"0490", X"03D2", X"0186", X"FED1", X"FF9B", X"03FB", X"04DE", X"061A", X"04A4", X"FF21", X"0105", X"043E", X"07E5", X"05F2", X"079D", X"024F", X"002A", X"FFB7", X"0231", X"04E7", X"02C0", X"0488", X"05B8", X"0358", X"02B4", X"0358", X"0484", X"0299", X"026A", X"0312", X"FF00", X"FE1E", X"FEBE", X"02AC", X"04DC", X"044B", X"0202", X"FF84", X"FE8A", X"FFE0", X"0017", X"029F", X"0583", X"FFF5", X"FFAE", X"00B2", X"01BE", X"027A", X"037D", X"026D", X"00F8", X"02EB", X"FF09", X"0015", X"00C1", X"02CC", X"FF8D", X"00F6", X"FD6E", X"FC96", X"FE7E", X"01D9", X"076A", X"05C4", X"0363", X"FF98", X"FFDE", X"FD90", X"FF8F", X"012E", X"019F", X"FC2B", X"FF7C", X"FFAA", X"FF22", X"FF2A", X"0220", X"00EA", X"FFA2", X"FD56", X"FC46", X"FCAF", X"FEA4", X"005B", X"01A0", X"FD96", X"FBC1", X"FC1E", X"004E", X"06E0", X"09E4", X"060E", X"034D", X"01C9", X"FF17", X"FE6D", X"FDE6", X"FEB3", X"FC3C", X"FD8A", X"FF5B", X"0100", X"FBD9", X"FDA8", X"0012", X"FE0F", X"FC8D", X"FB98", X"FB1F", X"FB2B", X"FC37", X"FC77", X"FEB5", X"FC25", X"FAB1", X"FC7B", X"0046", X"0610", X"061B", X"026C", X"00AF", X"00AC", X"FF98", X"FDA9", X"FEE5", X"FA55", X"FF10", X"FE11", X"00BF", X"005A", X"FDF4", X"FE73", X"FF2A", X"FD51", X"FDE8", X"FBBE", X"FBB5", X"F8BE", X"F8FE", X"F9D0", X"FCC7", X"FB89", X"F846", X"FCE5", X"02D5", X"061C", X"02B9", X"FFD0", X"FEFE", X"011E", X"FD64", X"FE10", X"FDDD", X"F8FA", X"FCA1", X"FFD9", X"008E", X"FF70", X"FD91", X"FFFA", X"00D3", X"FEFA", X"FFAC", X"FE22", X"FCAD", X"FB72", X"F86B", X"F92C", X"FCE1", X"F9FE", X"FAAD", X"FC72", X"0162", X"01B5", X"010E", X"FFE2", X"FF02", X"FDB7", X"FDFA", X"FE3D", X"0079", X"F8FA", X"FE09", X"01A0", X"0069", X"01A5", X"FFD1", X"FFF4", X"FF08", X"023C", X"019A", X"FEE0", X"FCDC", X"FD72", X"FCE2", X"FCE3", X"FC21", X"FD03", X"FBF0", X"FE3A", X"013C", X"FFAB", X"0029", X"FF4E", X"004C", X"FEEA", X"FF41", X"FCAC", X"FB0B", X"F675", X"FEC7", X"FDAF", X"00AD", X"013D", X"0205", X"003E", X"FFD9", X"0575", X"02DF", X"001B", X"FF6A", X"FCD8", X"FDF6", X"FC5E", X"FF81", X"FD05", X"FEC7", X"FD8C", X"FDC2", X"FEBC", X"FD2E", X"FF12", X"FE7E", X"FE83", X"FD81", X"FD95", X"FB89", X"F7B1", X"F9EE", X"FDB3", X"0093", X"0264", X"00A8", X"FFC6", X"FE31", X"0358", X"0194", X"FF70", X"FF59", X"FE78", X"FDB0", X"FB18", X"FE7E", X"FF52", X"FF6E", X"FEC9", X"FE2F", X"FDD6", X"FCBD", X"FCC3", X"FC5A", X"FDFF", X"FCFF", X"001D", X"FC38", X"FE0C", X"FA1D", X"010F", X"FFB8", X"FF98", X"02B1", X"FF97", X"FD2E", X"FFC1", X"013D", X"FF3A", X"004F", X"FF6B", X"FD9D", X"FCE3", X"FE79", X"00AA", X"FDBB", X"FE7E", X"FDD8", X"FC2D", X"FA61", X"FB43", X"FA8F", X"FDC8", X"0004", X"FEFF", X"FB44", X"FDD2", X"FC73", X"FFDC", X"FF22", X"FED0", X"0271", X"007A", X"FBB9", X"F99A", X"FFB0", X"01F2", X"0077", X"009A", X"018E", X"021C", X"03A8", X"0360", X"0250", X"FF7A", X"FE4F", X"FB70", X"F983", X"FA36", X"FA79", X"FEFD", X"046D", X"03C3", X"0148", X"FFC9", X"FF83", X"0078", X"00DD", X"0021", X"00C4", X"0402", X"0086", X"FCC3", X"FECF", X"0178", X"0336", X"0445", X"06A7", X"057B", X"0353", X"0512", X"0412", X"008E", X"00B5", X"FDE2", X"FFAA", X"FE94", X"00A4", X"026E", X"026F", X"0557", X"0384", X"0075", X"FE40", X"00F2", X"0068", X"FFFC", X"00C8", X"053A", X"039B", X"FF1F", X"0183", X"0217", X"054D", X"04C1", X"0549", X"0776", X"05B3", X"08FC", X"0887", X"074C", X"04E9", X"0301", X"02AC", X"04A5", X"025A", X"0114", X"02A5", X"05DB", X"0190", X"FC8A", X"FDBF", X"FFC7", X"0043", X"01AB", X"FFDD", X"03B9", X"054F", X"066A", X"0543", X"0516", X"069C", X"07EB", X"0982", X"08F1", X"077F", X"0A0A", X"0973", X"0B2D", X"0D3C", X"0C32", X"0A98", X"08D4", X"0664", X"03AA", X"037E", X"01EC", X"00C8", X"FF67", X"FED1", X"FEFF", X"FF15", X"FE9B", X"00D9", X"FFAE", X"FF80", X"0212", X"029A", X"01C7", X"0467", X"039B", X"035E", X"0418", X"06E2", X"072B", X"08F1", X"07B2", X"07F2", X"06FA", X"074D", X"05B3", X"04B4", X"03A1", X"01C3", X"0153", X"0217", X"00F0", X"FE8B", X"FE75", X"FFFF", X"0146", X"00E1", X"008B", X"FED3", X"005C", X"0083", X"01B4", X"01A8", X"0151", X"02FB", X"00F4", X"03C5", X"03CC", X"0416", X"01AF", X"FFB0", X"03E3", X"028D", X"01E1", X"0154", X"02D9", X"0168", X"00A3", X"FEC5", X"002B", X"FF29", X"FE6C"),
--        (X"00CF", X"FF99", X"00B0", X"01C4", X"011F", X"FECB", X"FEEB", X"FE82", X"0032", X"009E", X"FF9E", X"0003", X"043B", X"0209", X"0023", X"001D", X"0140", X"FF8A", X"FE60", X"0195", X"00E2", X"00B6", X"00A5", X"0024", X"003E", X"0021", X"FFEF", X"017C", X"FEC5", X"FFDF", X"0094", X"0008", X"00EF", X"0105", X"0564", X"051D", X"04C9", X"044B", X"074B", X"077F", X"074A", X"07DC", X"0103", X"028A", X"0223", X"053D", X"06B2", X"058D", X"0596", X"0443", X"03BB", X"02C8", X"0061", X"0089", X"FE9E", X"FFB3", X"FFC2", X"FE7F", X"00B1", X"0148", X"02A1", X"014C", X"0700", X"06F0", X"0A21", X"053D", X"0743", X"0816", X"0800", X"0525", X"04EF", X"0322", X"03B8", X"013F", X"00D6", X"023A", X"043C", X"03F9", X"0720", X"066F", X"0107", X"FE04", X"003E", X"FF7E", X"003F", X"002E", X"FF08", X"02C3", X"FF0A", X"04A6", X"02E6", X"0553", X"0584", X"0372", X"0389", X"05AA", X"0539", X"03D2", X"0259", X"0026", X"008D", X"00E7", X"0017", X"FFF7", X"0345", X"02F9", X"0329", X"035B", X"01B6", X"FD7A", X"01F0", X"FFBC", X"0146", X"FF77", X"FD6F", X"013D", X"0064", X"002A", X"FED0", X"0044", X"0163", X"00B6", X"00C0", X"001C", X"FFCC", X"0149", X"FF27", X"007C", X"FF1B", X"0028", X"FFC0", X"FE4E", X"00B6", X"00E5", X"0349", X"0330", X"FE02", X"FC8D", X"FE4B", X"0297", X"FFA6", X"FF1F", X"FD55", X"FB72", X"002D", X"FCC0", X"FF2F", X"FE4E", X"001B", X"FDD8", X"00CB", X"FE4E", X"FDF3", X"0178", X"0079", X"015B", X"FF0C", X"0069", X"0113", X"006D", X"FFDF", X"FE58", X"FF0A", X"FF78", X"FCC3", X"F8DC", X"FE42", X"0201", X"0048", X"0044", X"00FD", X"00BA", X"00AE", X"FD06", X"FFC8", X"FECE", X"FDEB", X"FBB9", X"FABE", X"FCA0", X"FFD2", X"FF3A", X"FE09", X"FDED", X"FCEC", X"FD7D", X"FE75", X"FDF3", X"FE2F", X"0005", X"FF4A", X"FCBA", X"F81A", X"F572", X"F787", X"FDC9", X"0021", X"0366", X"FEA4", X"FF50", X"019C", X"FEF2", X"FC6E", X"FD89", X"FA2B", X"FBA6", X"FAC1", X"FC80", X"FD1C", X"FBA3", X"FC8B", X"FB6D", X"FC6F", X"FF4F", X"FD70", X"FD22", X"FDE5", X"FE78", X"FDEF", X"FD1E", X"FB54", X"F66A", X"FB34", X"FD46", X"02F7", X"0256", X"00B6", X"02D7", X"026E", X"FF94", X"FDE5", X"FD8F", X"FBD9", X"FB95", X"FAFC", X"FAB2", X"FBF3", X"FC9B", X"FCA6", X"01BE", X"001F", X"FF80", X"FDEC", X"FC79", X"FD87", X"FDB3", X"FC79", X"FD4D", X"F998", X"F5F0", X"F99A", X"FDC1", X"017A", X"029F", X"044D", X"03CB", X"0381", X"FF84", X"FF2A", X"FF8E", X"FE0B", X"FCD4", X"FE8B", X"FCF1", X"FDB8", X"005F", X"0590", X"0447", X"010D", X"FDDE", X"FC3D", X"FDAE", X"FEC6", X"FF9D", X"FE4F", X"FF6F", X"FFAB", X"F7AD", X"FB92", X"FF76", X"01AA", X"0479", X"05B2", X"0563", X"008C", X"0124", X"FF96", X"FFD8", X"FF4C", X"FF0E", X"0120", X"01A3", X"012E", X"06CE", X"06C9", X"0197", X"FE1A", X"FC9D", X"FECF", X"FECF", X"0412", X"028B", X"028B", X"04FC", X"0210", X"FA98", X"FB6A", X"FE7B", X"027C", X"0608", X"0818", X"0424", X"0148", X"FF56", X"007A", X"021B", X"029F", X"044D", X"0480", X"03D5", X"0643", X"098F", X"01BA", X"F8C9", X"F95A", X"FCEE", X"FF85", X"0129", X"03C5", X"03AA", X"0431", X"0581", X"04A8", X"FB38", X"F77F", X"FE82", X"0158", X"048B", X"07D6", X"008D", X"FF9D", X"01D0", X"03F8", X"066B", X"0566", X"0779", X"058D", X"05F5", X"05AA", X"025E", X"FC75", X"F9EF", X"FCC7", X"FEBB", X"005D", X"007E", X"014F", X"01D0", X"03BE", X"060C", X"0422", X"FC59", X"F8B6", X"FE3E", X"0032", X"017C", X"0878", X"FFD6", X"FFE4", X"046C", X"0787", X"0649", X"05A5", X"0498", X"0467", X"002B", X"0222", X"FAA0", X"F8C7", X"FBEA", X"FE6F", X"FE56", X"00CB", X"FFE0", X"003A", X"0145", X"0041", X"0677", X"036E", X"FC81", X"F639", X"FAA2", X"002A", X"00E7", X"0417", X"FD54", X"FC77", X"039B", X"0482", X"0525", X"0381", X"02EC", X"0094", X"FF9B", X"FD58", X"FA3A", X"FAA8", X"FDEA", X"FC51", X"FC08", X"FEF0", X"0077", X"FF98", X"00C5", X"00E6", X"036F", X"00F6", X"F945", X"F825", X"FCE1", X"0040", X"FFE4", X"021E", X"F9EE", X"FBC5", X"00A7", X"0199", X"03D7", X"03B6", X"0168", X"00FA", X"0163", X"FB27", X"F9EB", X"FAA2", X"FBFF", X"FA8A", X"FD72", X"FF73", X"FF8C", X"0118", X"FEC5", X"0080", X"0267", X"00B2", X"FC08", X"F725", X"FBD8", X"00CB", X"017B", X"FE74", X"F935", X"FBA9", X"0051", X"FF3F", X"03DD", X"035E", X"0254", X"0171", X"019D", X"F90B", X"F980", X"FA74", X"FA56", X"FA3A", X"FBCE", X"FE2B", X"0011", X"FF3B", X"FF0C", X"FDE1", X"0092", X"0195", X"FB70", X"F66B", X"FB40", X"FFB8", X"0000", X"FC35", X"F8E4", X"FBA4", X"FDBA", X"FD3E", X"01F7", X"022A", X"03A9", X"038B", X"02DF", X"FE01", X"FAA5", X"FA7B", X"F9A0", X"FAB8", X"FF4A", X"FE9A", X"FF3A", X"00D2", X"FF1A", X"00DA", X"01C8", X"FF6B", X"FE7D", X"FA55", X"FF23", X"0193", X"0061", X"FE0B", X"F9A1", X"FC34", X"FB61", X"FB77", X"FF24", X"042D", X"02BA", X"05A2", X"0459", X"04D2", X"FEE2", X"FCEC", X"FC80", X"FDBD", X"00E2", X"FEE8", X"FF1A", X"00D5", X"FEEA", X"00EF", X"FFDC", X"FCD5", X"0095", X"FCCC", X"FDFA", X"FFA5", X"032A", X"FEB3", X"F8DB", X"FB40", X"FB82", X"FB3B", X"FEDB", X"00C0", X"03D5", X"0518", X"0903", X"08B0", X"0473", X"0001", X"FFBC", X"FFCF", X"FF9F", X"FFD9", X"013D", X"0051", X"00C7", X"00E6", X"FFBF", X"FDB7", X"FCD5", X"FC3E", X"FD2C", X"0033", X"0254", X"FD7E", X"F70F", X"FCF3", X"FDC8", X"FB46", X"FD08", X"FEA7", X"0044", X"01B0", X"04A8", X"0741", X"0678", X"049C", X"0154", X"FFA7", X"FFB2", X"FF43", X"FEF6", X"000A", X"FE40", X"FD82", X"FD9F", X"FD2F", X"FC71", X"00F7", X"002C", X"FF14", X"0035", X"FD5E", X"F88B", X"FB2B", X"FCD1", X"FB65", X"FBED", X"FCDA", X"FE6C", X"0128", X"01FC", X"03AA", X"0424", X"0473", X"024B", X"00D8", X"0030", X"FFA5", X"FDF4", X"0000", X"FEB2", X"0087", X"FD6B", X"FDD2", X"FE46", X"02DE", X"FFE8", X"002A", X"FF55", X"FED9", X"FB56", X"F85B", X"FBD4", X"FD27", X"FC78", X"FF6E", X"0017", X"FF9D", X"0192", X"04EB", X"0454", X"02BA", X"02FC", X"0192", X"01AB", X"FFE9", X"FFE5", X"FFBF", X"FF50", X"FF75", X"FC1B", X"F966", X"FC88", X"049C", X"0090", X"FF29", X"FFC3", X"02B9", X"FC87", X"FB85", X"FD89", X"FE6D", X"FF2D", X"0018", X"0215", X"01EB", X"0239", X"031A", X"0145", X"03C6", X"036D", X"FF9D", X"0177", X"FE1B", X"FCA4", X"FDA1", X"FDBE", X"FBD7", X"F9B2", X"F95D", X"FC52", X"01AB", X"FE5A", X"FF02", X"FE87", X"01ED", X"01E6", X"015F", X"000A", X"FD57", X"FD02", X"FDE6", X"FEC8", X"FEB1", X"FF95", X"FF6A", X"FEEF", X"0021", X"FE57", X"FEF5", X"FF42", X"FCE9", X"F9C7", X"F9DD", X"FB64", X"FBD3", X"F880", X"FC10", X"FEA3", X"0092", X"FF3E", X"FFC2", X"002A", X"FE09", X"0321", X"0273", X"FF0D", X"FC40", X"FC03", X"FE13", X"FA92", X"FAD4", X"FC20", X"FB80", X"FA45", X"F904", X"FA89", X"FCEE", X"FE5C", X"FE38", X"FE5B", X"FE2E", X"FF27", X"FF41", X"FBF5", X"0078", X"FFD0", X"005A", X"FF4F", X"0001", X"004B", X"0000", X"0066", X"FD0D", X"FE15", X"FFEC", X"00BB", X"02DF", X"FF83", X"FFA1", X"023A", X"0016", X"00EB", X"FEF2", X"0182", X"04E2", X"05A0", X"0245", X"0571", X"019D", X"02FF", X"0566", X"FFDD", X"FFA9", X"01DE", X"00D2", X"0144", X"00EA", X"FFEF", X"00C4", X"FEDD", X"0418", X"01DD", X"0215", X"FF62", X"036E", X"0426", X"022D", X"01D5", X"FF93", X"05A7", X"01DD", X"014C", X"058E", X"04DF", X"02FD", X"051E", X"02BD", X"03C9", X"0420", X"02E3", X"00EA", X"009C", X"FFAC", X"FF40"),
--        (X"FF0D", X"FFB5", X"FF27", X"FFC1", X"016B", X"003F", X"FFA1", X"FFE3", X"FFA0", X"00DA", X"00AA", X"FFC9", X"0107", X"FFDD", X"FF10", X"012E", X"000C", X"0179", X"FDF5", X"0108", X"003E", X"FE8E", X"FF67", X"008A", X"0058", X"006C", X"FF73", X"FFE5", X"FFFD", X"00C3", X"002D", X"FF83", X"003F", X"0044", X"006E", X"0016", X"FEE9", X"FD96", X"FE4F", X"FDD3", X"FE89", X"FEB7", X"002F", X"01C9", X"FE16", X"FCC1", X"FF5E", X"FFCE", X"FD80", X"0049", X"0108", X"FEDB", X"FF8D", X"FEAA", X"FFA9", X"FF77", X"0130", X"00A8", X"FF84", X"0069", X"001A", X"0158", X"FDCE", X"FF22", X"FC0D", X"F886", X"FA14", X"FC6E", X"003A", X"FD8D", X"FEB3", X"FD93", X"FFF5", X"FECB", X"FF50", X"001D", X"FE6B", X"FC87", X"FE20", X"FD91", X"FC3C", X"FF86", X"0074", X"00A1", X"FF53", X"000D", X"027C", X"0312", X"0235", X"010D", X"FF34", X"000D", X"0172", X"FE89", X"FE66", X"FD33", X"FFC7", X"FF45", X"FDDA", X"FEF3", X"FED3", X"FF1D", X"0084", X"FF43", X"0224", X"FED9", X"FE27", X"FF0A", X"FD13", X"FEA7", X"FEA0", X"000E", X"FE15", X"00C5", X"0317", X"038E", X"0430", X"025D", X"019C", X"027B", X"0286", X"FE62", X"FE7D", X"FEBF", X"FF97", X"0259", X"018A", X"01E8", X"0138", X"00C3", X"01AF", X"0177", X"00C0", X"014A", X"FEC8", X"FD77", X"FDB6", X"FD22", X"FE32", X"FDBB", X"FEED", X"FFDF", X"0127", X"01E5", X"0257", X"0392", X"017A", X"FF08", X"FD5B", X"FD6D", X"FCE8", X"FC5F", X"FE13", X"FF4A", X"FF83", X"0142", X"0202", X"017A", X"00F5", X"0190", X"0294", X"0022", X"FFB5", X"FF9B", X"FCDD", X"FEEC", X"0021", X"FE23", X"FF62", X"00F6", X"0107", X"0156", X"0251", X"019A", X"0045", X"FF03", X"FD04", X"FD6F", X"FD29", X"FD2A", X"FED3", X"FF48", X"FE4B", X"FF0D", X"FE66", X"0042", X"01BB", X"0161", X"01C6", X"0010", X"FEC9", X"FF00", X"02AB", X"0070", X"0219", X"FEAB", X"0010", X"00EC", X"FD87", X"FFAB", X"024C", X"0219", X"FF62", X"FF72", X"FF07", X"FD28", X"FD8D", X"FDAA", X"FDB6", X"FEE5", X"0019", X"FDE0", X"FF24", X"FF5C", X"0038", X"00B4", X"001A", X"FD34", X"FE21", X"FEE8", X"FF28", X"041D", X"023D", X"FF52", X"FEDB", X"FC40", X"FC9D", X"004C", X"01DF", X"FFCB", X"FDA3", X"FD51", X"FE2B", X"0013", X"FF9C", X"FEB7", X"FFFE", X"FE22", X"FF7B", X"FF1F", X"FEFC", X"FF7D", X"FF38", X"FEA4", X"FDF2", X"FFFA", X"013E", X"0013", X"034C", X"0916", X"0578", X"018B", X"FD49", X"FC53", X"FD41", X"FE33", X"FF14", X"FDA6", X"FCFD", X"FF24", X"FEDD", X"018F", X"013A", X"0267", X"01A4", X"0187", X"FE18", X"0084", X"FEDE", X"0124", X"FF26", X"FF5A", X"FF0A", X"0053", X"017B", X"013B", X"0423", X"07D0", X"05B0", X"FE9E", X"FFF0", X"FE20", X"FC68", X"0099", X"FFFA", X"FB5B", X"FB78", X"FD9D", X"FF2F", X"FFE8", X"0024", X"0230", X"025F", X"02F4", X"03FB", X"03F1", X"0127", X"01FB", X"FE71", X"FE7D", X"FE6F", X"FE52", X"0275", X"01E2", X"06D4", X"0A22", X"038F", X"FEF9", X"0009", X"FBA1", X"FB6A", X"FF19", X"FD54", X"F8A0", X"F7A2", X"F9E2", X"FC76", X"FD6A", X"FF19", X"01AB", X"0547", X"05F0", X"054D", X"0515", X"04A6", X"03B0", X"020C", X"FF48", X"FE4D", X"FB8E", X"FA1C", X"FF4D", X"0189", X"0870", X"0650", X"FFA7", X"FEDC", X"FB76", X"F928", X"FBAF", X"FC7A", X"F7D2", X"F876", X"F8C6", X"FA5F", X"FBFD", X"00B2", X"02BB", X"0627", X"0579", X"0636", X"0444", X"055C", X"0329", X"01D6", X"FF04", X"FD88", X"F7F6", X"F6D3", X"F611", X"F7F2", X"FF28", X"0178", X"FE68", X"00B8", X"FCAF", X"F9BF", X"FC87", X"FE3B", X"F8EB", X"F73F", X"F7CD", X"F9C6", X"FB7B", X"FA73", X"0140", X"040F", X"0676", X"04DE", X"0419", X"0422", X"00A7", X"FFF6", X"00F9", X"FC24", X"F82E", X"F6C0", X"F534", X"F589", X"F995", X"FB82", X"FCF5", X"005A", X"0177", X"FDD8", X"FFA1", X"FDD8", X"F97D", X"F4E3", X"F52F", X"F6B0", X"F788", X"F921", X"FC32", X"03AE", X"0620", X"0571", X"03DE", X"007F", X"FFA6", X"FE14", X"FF7A", X"FE6E", X"FDCF", X"FAE5", X"F919", X"F6EB", X"FB60", X"FD03", X"FF90", X"0122", X"011C", X"000E", X"FE31", X"FEB6", X"FAC6", X"F824", X"F4F9", X"F53F", X"F40D", X"F4FF", X"FADF", X"01F4", X"03B5", X"01F9", X"0178", X"FDEF", X"FE57", X"FF86", X"0140", X"0127", X"0126", X"0120", X"FC2A", X"F806", X"F90D", X"FC0E", X"FEBF", X"FEED", X"02DF", X"00E8", X"01C4", X"035D", X"00F6", X"FE2C", X"F869", X"F4B0", X"F377", X"F242", X"F645", X"FB9A", X"0084", X"FFCE", X"FE14", X"FE1C", X"FCDC", X"FF94", X"0287", X"0233", X"01EA", X"FFFF", X"FC6B", X"F94D", X"F62A", X"FCAC", X"FDA6", X"0002", X"029F", X"FFC9", X"03E7", X"060F", X"03F5", X"030F", X"FF80", X"FA55", X"F4DE", X"F5AE", X"F2F0", X"F736", X"F9C3", X"FEB6", X"FEC3", X"FFB7", X"008B", X"FFB5", X"02F7", X"03BA", X"0452", X"0090", X"FC3A", X"F754", X"F719", X"FC46", X"FB85", X"FE93", X"022A", X"FF20", X"0632", X"059F", X"03A9", X"052A", X"00CE", X"003D", X"FDC3", X"F99A", X"F843", X"F85F", X"F958", X"FDFA", X"0076", X"00B7", X"0181", X"0238", X"00B5", X"02F3", X"01C7", X"FE02", X"F9F9", X"F722", X"FB54", X"FE0D", X"01AB", X"0070", X"FDB0", X"FE68", X"0468", X"035D", X"034D", X"02DB", X"0294", X"0461", X"02FD", X"00EA", X"FDDA", X"FBF9", X"FDB8", X"FF18", X"0056", X"01D3", X"022D", X"01FB", X"01D6", X"016C", X"FFFB", X"FD99", X"FA34", X"FB6B", X"FE27", X"FF78", X"007B", X"FFA4", X"0039", X"FD99", X"0051", X"01A8", X"0206", X"04C8", X"0251", X"0480", X"01C1", X"0263", X"005C", X"FDE6", X"FE33", X"FFFC", X"FF85", X"010A", X"0265", X"0289", X"FFB2", X"FF7E", X"FF8E", X"FC29", X"FB01", X"FAA5", X"FE99", X"FF3D", X"0136", X"0053", X"0192", X"000D", X"0022", X"01BF", X"021E", X"0322", X"03FF", X"01F8", X"03B4", X"0342", X"FFAC", X"FED2", X"FCAB", X"FEEC", X"0039", X"FEB6", X"FF01", X"0055", X"FFC3", X"0145", X"FD7F", X"F8F2", X"F6B9", X"FBA9", X"FA15", X"FFA9", X"FDCD", X"0122", X"01EA", X"00B4", X"003B", X"02B7", X"FFAC", X"00C0", X"FE10", X"000B", X"FF78", X"0158", X"FFC4", X"FDEE", X"FE32", X"FE67", X"FEA6", X"0027", X"025F", X"0029", X"FF82", X"FED3", X"FB3B", X"F795", X"F9D3", X"F8DB", X"FA68", X"027D", X"010E", X"FFAB", X"0034", X"02B1", X"0459", X"0465", X"03A2", X"00B4", X"0016", X"FE2C", X"FFE9", X"FFBC", X"011F", X"0116", X"0123", X"FFD8", X"010C", X"FF7C", X"FFB3", X"FDD2", X"FDC0", X"FC20", X"F7BD", X"F75B", X"F9AE", X"FFA4", X"0039", X"03EA", X"005C", X"FFF8", X"FFF7", X"FF4C", X"042D", X"0236", X"FFFD", X"01E4", X"025F", X"02CE", X"02EB", X"0239", X"01C3", X"FFB8", X"FF12", X"FF8F", X"FE1F", X"FEFD", X"FEA4", X"F955", X"FB02", X"FB9F", X"FB49", X"FB5A", X"FE2A", X"FC67", X"002E", X"0104", X"FF7C", X"0037", X"00EA", X"0076", X"FE2D", X"FE36", X"FD43", X"000C", X"01A3", X"0413", X"01DC", X"013A", X"FF4A", X"FEE7", X"FF33", X"FB69", X"F9E6", X"F91A", X"F85E", X"F9DC", X"FCA1", X"FF14", X"FE6D", X"FFA6", X"FC3A", X"FF36", X"0041", X"FED0", X"FFBB", X"00EB", X"FFFB", X"00CE", X"01B1", X"014E", X"FD1F", X"FD6D", X"FCF7", X"FC44", X"FCBF", X"FC1C", X"FC57", X"FAF2", X"FA07", X"F9CF", X"FBED", X"FC54", X"FACE", X"FB37", X"FBAD", X"FEE2", X"0058", X"FF79", X"FE17", X"FF86", X"FF5C", X"FEEE", X"0024", X"0057", X"FFA6", X"FF43", X"FFB5", X"FF05", X"000C", X"FF1C", X"FBFA", X"FB27", X"FDB1", X"FAB3", X"FAA4", X"FA33", X"F8AE", X"FD5A", X"FEE0", X"FB34", X"FACE", X"FCD5", X"F98C", X"FC49", X"FD10", X"FF6B", X"FEC7", X"005F", X"00D1", X"FF7C", X"0083"),
--        (X"FFAE", X"FFB5", X"FEFB", X"00AA", X"00A2", X"FFF5", X"005C", X"001B", X"FF9C", X"01C9", X"0048", X"0001", X"00EB", X"0071", X"00A2", X"FDF8", X"01C2", X"FEA8", X"FF88", X"0192", X"FFEB", X"0210", X"FF58", X"0108", X"FF06", X"FFAC", X"00CC", X"FF21", X"FF74", X"FF32", X"FF39", X"000D", X"001F", X"FF84", X"03C5", X"036E", X"0001", X"FD12", X"FF62", X"FDC8", X"FE66", X"FE9D", X"0100", X"0192", X"007E", X"FFBF", X"FEC7", X"01A0", X"004E", X"0218", X"02F5", X"0392", X"FF5A", X"FF15", X"FECA", X"0003", X"00C5", X"FF54", X"0122", X"00BD", X"FFAA", X"00A3", X"0371", X"04A3", X"01FF", X"02E3", X"00AE", X"00AB", X"018F", X"FFBB", X"FE61", X"0141", X"0087", X"0258", X"026A", X"01A7", X"007E", X"FFB4", X"00CE", X"022B", X"FFB9", X"0111", X"FF94", X"FF18", X"FEB5", X"006C", X"000F", X"042D", X"0331", X"034F", X"01E5", X"00E7", X"FFEE", X"0040", X"0248", X"FFFD", X"015F", X"01A5", X"0109", X"0349", X"042D", X"015B", X"01DA", X"01CB", X"01DD", X"01DE", X"00A4", X"0030", X"00BA", X"0048", X"0014", X"FF23", X"00B6", X"0058", X"009C", X"00A4", X"FDAA", X"0220", X"0065", X"FDF4", X"009A", X"0031", X"01CB", X"0135", X"01DC", X"FF89", X"0450", X"0363", X"0436", X"01F3", X"0256", X"0108", X"FDF9", X"FE50", X"FD0C", X"FE0D", X"FF95", X"0374", X"0224", X"00CA", X"FFCB", X"FEA9", X"0127", X"026C", X"FFA1", X"004B", X"003B", X"012C", X"0079", X"00B9", X"FED6", X"FCCD", X"FD86", X"FE71", X"FEB3", X"FEB6", X"014A", X"014C", X"027E", X"015E", X"023D", X"00B7", X"0023", X"01A1", X"033C", X"0719", X"054C", X"029B", X"FE63", X"00F0", X"FE75", X"011F", X"0112", X"01BF", X"FFB5", X"0187", X"005F", X"FF7D", X"FE5C", X"FE80", X"FE39", X"FCF7", X"FE0F", X"001C", X"0014", X"00A7", X"FFC0", X"FFA1", X"0069", X"015C", X"FFD0", X"0292", X"0650", X"09D4", X"096E", X"035E", X"012C", X"022B", X"FEBE", X"FE70", X"02A5", X"013A", X"0090", X"01EE", X"00D1", X"FF0F", X"FF0A", X"FE00", X"FC5A", X"FF61", X"FEA1", X"FE0D", X"002D", X"FE83", X"FF1C", X"FF78", X"0068", X"0041", X"00A0", X"004D", X"04A4", X"0806", X"053A", X"0280", X"FFA5", X"FF8A", X"FCDC", X"FE61", X"01D3", X"0301", X"00D5", X"028D", X"FFFE", X"0088", X"0032", X"00AA", X"0146", X"01AD", X"00E0", X"FF90", X"0026", X"0035", X"FE35", X"00BB", X"FFCB", X"FFF0", X"0045", X"01A7", X"0310", X"093F", X"0656", X"04B0", X"0084", X"FDCC", X"FEFB", X"019C", X"019B", X"01F9", X"023B", X"0023", X"FEBB", X"FE33", X"007B", X"FFB7", X"0116", X"005E", X"0065", X"FFF2", X"FD63", X"FE0D", X"FE0D", X"FF3C", X"FF92", X"0034", X"017F", X"FEAD", X"039F", X"0BBE", X"0A00", X"021C", X"00A0", X"FCD3", X"FE1F", X"0341", X"01CE", X"FF43", X"00C1", X"0055", X"FEA7", X"FF41", X"FDE4", X"FD46", X"FEC5", X"0123", X"0281", X"00B9", X"FD08", X"FAAB", X"FE26", X"FDAD", X"FCB5", X"FE79", X"FE0F", X"FE75", X"0500", X"0AED", X"08DA", X"0134", X"FF37", X"FE06", X"0072", X"0112", X"0116", X"00C2", X"FEE5", X"FF65", X"FE08", X"FBA0", X"FBFB", X"FA2A", X"FD66", X"0317", X"06B3", X"0201", X"FB34", X"F71C", X"FBEA", X"FE29", X"FBA6", X"FB04", X"FB77", X"FDB9", X"0251", X"0D2B", X"0849", X"012F", X"010F", X"FF34", X"FE2F", X"00D2", X"FE72", X"FE6A", X"FB46", X"FC25", X"FB23", X"FAF3", X"F9CB", X"FA5B", X"0108", X"06B4", X"0751", X"01E0", X"FB3E", X"F7FA", X"FC9A", X"FC93", X"FD74", X"FCE5", X"F971", X"FA3B", X"FC29", X"0927", X"0659", X"0174", X"00FF", X"FDF7", X"FF19", X"0046", X"FABE", X"F8D2", X"FB4F", X"F9E2", X"FA90", X"FC02", X"FA73", X"FD4A", X"04EB", X"0A38", X"06D0", X"0235", X"FC8D", X"FBC8", X"FEC3", X"FFFD", X"0013", X"FBE4", X"F896", X"FBB3", X"FBF6", X"0536", X"0743", X"032C", X"00C1", X"FF81", X"FF3F", X"FDBD", X"F9AD", X"F88A", X"FCBC", X"FB40", X"FBF4", X"FC97", X"FC96", X"0294", X"0704", X"095D", X"0700", X"034B", X"FBE7", X"FD36", X"FFB6", X"FEAC", X"FF5D", X"FCAB", X"FB22", X"FB15", X"FD6D", X"05CE", X"0460", X"0138", X"0215", X"FF0F", X"0162", X"00C4", X"FBB1", X"FB87", X"FD9C", X"FC5F", X"FC5B", X"FD98", X"0000", X"022C", X"098F", X"0A5B", X"075A", X"02D0", X"FEDE", X"FD17", X"FEDD", X"FFCA", X"FF18", X"0073", X"FAF9", X"FB2F", X"0244", X"06F4", X"02C9", X"00C0", X"FE4A", X"004B", X"020D", X"05F4", X"0286", X"FF17", X"FFF0", X"FB8C", X"FCC9", X"FEC8", X"00FD", X"05D3", X"0852", X"09A4", X"0816", X"01A6", X"FD75", X"FD6B", X"FE1E", X"015B", X"FFD7", X"002A", X"0163", X"015B", X"064F", X"070C", X"050E", X"0333", X"FF03", X"FF2E", X"0220", X"07B1", X"0486", X"00A2", X"0063", X"FEBC", X"FEED", X"FF06", X"0097", X"0524", X"0691", X"064A", X"01BB", X"FDD2", X"FFB8", X"FF0B", X"FEC9", X"01AA", X"FF1A", X"0188", X"FF3C", X"0470", X"0694", X"06C6", X"042B", X"0018", X"FD8E", X"008A", X"012C", X"0702", X"0365", X"0361", X"01E8", X"009D", X"FF57", X"00DB", X"FFFD", X"030B", X"0527", X"0432", X"00F7", X"FE39", X"FF14", X"011B", X"00BB", X"FE75", X"0003", X"0050", X"0337", X"05D8", X"0610", X"069F", X"02F0", X"0347", X"FF75", X"0035", X"FE74", X"03E4", X"0099", X"0268", X"01BD", X"00D4", X"02D0", X"0210", X"01EF", X"0224", X"0358", X"02D9", X"0136", X"01D0", X"018A", X"013C", X"01C9", X"004A", X"022E", X"028A", X"02C7", X"05C4", X"0305", X"0525", X"040F", X"FFCC", X"FF12", X"FD50", X"FF09", X"0306", X"01AE", X"0101", X"02F9", X"04A5", X"0495", X"0382", X"029D", X"0047", X"FFAF", X"007E", X"016C", X"01AB", X"01B9", X"004A", X"0212", X"006B", X"03C5", X"04CD", X"03D7", X"0528", X"01CA", X"FFDF", X"0114", X"FEAA", X"0121", X"0067", X"0535", X"0454", X"01A9", X"FED7", X"0068", X"01B8", X"044C", X"0136", X"00CE", X"FF15", X"FFEE", X"013C", X"021D", X"01D3", X"00D2", X"023B", X"01B2", X"02B4", X"02C5", X"00FB", X"030F", X"0492", X"00C3", X"01AD", X"014D", X"002E", X"0016", X"003B", X"05E0", X"0548", X"04ED", X"0108", X"0249", X"02A6", X"00F2", X"023E", X"FF88", X"005C", X"FF2D", X"FE8B", X"012D", X"FFCA", X"FFA3", X"018C", X"027D", X"022D", X"0377", X"00D0", X"FF23", X"FFA0", X"0069", X"00D6", X"00DD", X"FF79", X"FF72", X"018A", X"04FD", X"05C5", X"073C", X"028C", X"022A", X"0094", X"0165", X"01A9", X"FEBF", X"FF77", X"014D", X"0025", X"003B", X"01E1", X"034F", X"0111", X"0114", X"0316", X"0071", X"FED5", X"0073", X"FEFA", X"FFCD", X"000B", X"03B9", X"FFBA", X"FFCB", X"003D", X"0271", X"0371", X"0028", X"FCDA", X"FF99", X"FF6C", X"01A2", X"FFD0", X"FF4E", X"00D9", X"01C3", X"02F0", X"03B3", X"0292", X"01D0", X"01D2", X"0208", X"0100", X"FCCD", X"FC5A", X"FCE8", X"FF3A", X"02CB", X"0041", X"010F", X"0069", X"0062", X"FEB2", X"0245", X"FFB2", X"FC1D", X"FC5D", X"FD11", X"FC9A", X"FDE1", X"013D", X"0099", X"0222", X"01F1", X"02DB", X"01E3", X"021D", X"026B", X"013A", X"FFC7", X"FFF6", X"FD43", X"FB54", X"FE71", X"01B5", X"0426", X"FEF1", X"01AD", X"FF0F", X"FFDE", X"00C4", X"FF85", X"FD8D", X"F8D2", X"F9CE", X"F817", X"FB5A", X"F86E", X"FAB4", X"FBA8", X"FC19", X"FB49", X"FA5B", X"F936", X"FA51", X"FA81", X"FB99", X"FBA9", X"FD3D", X"F8A3", X"F8A3", X"FB1F", X"FCB0", X"FE46", X"FF26", X"002C", X"FED6", X"FFB0", X"002B", X"FFA6", X"001D", X"FFFC", X"FF08", X"FCEF", X"FD01", X"FD1E", X"FC48", X"FCEF", X"FF5B", X"FDF6", X"FCCD", X"F9FC", X"FA47", X"FC55", X"FD2A", X"FCE7", X"FBC9", X"FC63", X"FC2B", X"FD9E", X"003E", X"01B6", X"FFC8", X"FFDF", X"FF2D"),
--        (X"001F", X"0143", X"0067", X"004B", X"0026", X"0080", X"003F", X"0215", X"FF42", X"001C", X"FF53", X"0035", X"FF54", X"FE98", X"FE67", X"FF06", X"FE9C", X"FF7D", X"FE1A", X"0034", X"FF46", X"000C", X"FF30", X"0038", X"0123", X"00E4", X"FF92", X"00AB", X"FFBE", X"FF47", X"0086", X"FF6F", X"FF97", X"FFE3", X"00CB", X"0261", X"019D", X"042C", X"03B6", X"0630", X"05A2", X"05E5", X"FFA3", X"FE4F", X"0117", X"0486", X"045A", X"04CE", X"0471", X"03C9", X"0359", X"0169", X"FEBE", X"FE8D", X"FFE6", X"0018", X"0038", X"0113", X"0096", X"02B8", X"0216", X"0143", X"0252", X"018C", X"038D", X"02AA", X"03EA", X"0598", X"03B9", X"03EA", X"0209", X"033C", X"005E", X"00E2", X"017F", X"060C", X"058E", X"066A", X"06D8", X"0509", X"0399", X"0094", X"FF76", X"FF84", X"0122", X"FFE6", X"FDC0", X"03AB", X"0184", X"0444", X"03B6", X"049B", X"01EC", X"005D", X"03A1", X"0520", X"04AE", X"021D", X"0409", X"01D1", X"014A", X"0199", X"0340", X"0569", X"04B7", X"05CB", X"043E", X"03BF", X"0513", X"FFFD", X"FFB9", X"0223", X"0047", X"0001", X"0074", X"0466", X"032B", X"0275", X"0206", X"02FE", X"0327", X"FF59", X"021F", X"0117", X"FFAD", X"FEDC", X"FDA8", X"FE16", X"FD51", X"FF5F", X"01F9", X"030C", X"035F", X"0612", X"0723", X"04BF", X"00E7", X"FF68", X"FF68", X"FF2F", X"FF9A", X"FF19", X"01DE", X"02B6", X"037A", X"0471", X"031E", X"0224", X"0354", X"030D", X"00B1", X"FECE", X"FEE4", X"FF4A", X"FFD0", X"FFBF", X"FFD5", X"FFD7", X"001E", X"01A4", X"0058", X"01CE", X"0109", X"0420", X"00D3", X"FECF", X"FEEC", X"FEC3", X"FF15", X"0093", X"0462", X"04EA", X"041B", X"0515", X"02B5", X"0263", X"01EB", X"0061", X"0208", X"0049", X"017F", X"012C", X"0203", X"0066", X"01B0", X"0206", X"029D", X"018F", X"008C", X"0091", X"0179", X"006C", X"FFBC", X"FF73", X"0111", X"FF3B", X"016D", X"0290", X"FFEA", X"0444", X"0483", X"0311", X"002D", X"FFD9", X"FF69", X"FFF3", X"FEAD", X"FF60", X"0037", X"0203", X"03A0", X"03C4", X"03ED", X"03B1", X"028D", X"FFBB", X"000F", X"FD78", X"FD0E", X"FAD2", X"FBD3", X"FE23", X"FFA8", X"FF45", X"0183", X"0123", X"000B", X"02D9", X"0276", X"0030", X"FFA0", X"FEB4", X"FF94", X"FF49", X"FD71", X"FF54", X"FFA1", X"FF08", X"01BD", X"0093", X"01F5", X"FF5C", X"FF8A", X"FDAD", X"FCE0", X"FCD8", X"FA62", X"F8DC", X"F9A4", X"FC7C", X"FBC2", X"FDF9", X"FF55", X"01F2", X"01F3", X"022C", X"0037", X"FD78", X"FD75", X"FF3F", X"FF15", X"FD2D", X"FDFA", X"FC3E", X"FF0F", X"FF1F", X"00D6", X"FF93", X"FE92", X"FEB0", X"FEFD", X"FF9A", X"FEB5", X"FC86", X"FC80", X"F886", X"FAF8", X"FA26", X"FE7D", X"0046", X"FDB1", X"005E", X"012C", X"03AE", X"FF3B", X"FE89", X"FCC8", X"FCE9", X"FCA7", X"FDA3", X"FC8D", X"FDF8", X"FE16", X"FE63", X"FC1F", X"FAC9", X"FC8C", X"00A1", X"FF42", X"FEBB", X"FFB6", X"FDB9", X"FC1E", X"FA39", X"FBC2", X"FF3E", X"FF3E", X"FF4B", X"FE9A", X"FF8A", X"05C6", X"0534", X"015B", X"FD5C", X"FE88", X"FDBD", X"FEB4", X"FCA8", X"00F4", X"0187", X"01A0", X"FEDE", X"FBA4", X"FC46", X"0221", X"03C7", X"0461", X"0142", X"030B", X"00B7", X"FE68", X"FEBD", X"FB95", X"FA96", X"FB0C", X"FFD4", X"FF0F", X"FF32", X"0348", X"0372", X"0023", X"0145", X"030E", X"0078", X"00BD", X"00C1", X"0581", X"04CD", X"01A3", X"005C", X"FD5B", X"FEAF", X"03C5", X"05D8", X"05C0", X"00F5", X"0221", X"02A4", X"0332", X"02D5", X"FF7B", X"F9C6", X"FA11", X"FED5", X"FDFD", X"0023", X"0028", X"0494", X"044F", X"060C", X"0840", X"087D", X"03C8", X"01F4", X"035B", X"0240", X"0126", X"FEB1", X"FD0C", X"FD79", X"0236", X"047C", X"029C", X"0369", X"0217", X"0277", X"0559", X"02CD", X"0007", X"F7D2", X"F8EB", X"FC26", X"0064", X"0343", X"0324", X"05F5", X"0901", X"0B56", X"0752", X"07AB", X"01A7", X"02E6", X"FF46", X"0084", X"FED5", X"FB9F", X"FC78", X"FD65", X"01EE", X"0282", X"0126", X"03E1", X"0461", X"0484", X"051F", X"0433", X"00A0", X"FA02", X"F7AD", X"FD9B", X"FF9B", X"02ED", X"00F6", X"02E9", X"05B4", X"0895", X"0626", X"04E2", X"02D6", X"00FD", X"00E4", X"0009", X"FD43", X"FB33", X"FBB0", X"FDCB", X"FEA0", X"00CA", X"01B8", X"043A", X"07CD", X"04BB", X"0462", X"027C", X"FCC6", X"F8A9", X"F9B5", X"FDDB", X"0042", X"01A1", X"001E", X"006C", X"057B", X"0554", X"FE9D", X"00C8", X"023B", X"FFD2", X"FF62", X"002C", X"FCF8", X"FC57", X"FA5C", X"FB4B", X"FC0F", X"018E", X"0315", X"061F", X"0649", X"026A", X"0355", X"0095", X"FD0E", X"F859", X"F75F", X"FE01", X"0009", X"0234", X"0171", X"FFF7", X"02A9", X"01DC", X"FEBD", X"FF57", X"FE4A", X"FDCD", X"FDBD", X"FE38", X"FCD1", X"FAEA", X"F8E1", X"FBDC", X"0033", X"048D", X"065A", X"05F5", X"FF26", X"0118", X"00F4", X"FDFD", X"FBAE", X"F8F3", X"FA4B", X"FD24", X"FE83", X"011F", X"01AC", X"0103", X"0447", X"FF92", X"FBE0", X"FC6A", X"FCCE", X"FEFA", X"FC30", X"FE68", X"FAAD", X"F74B", X"FAB0", X"003C", X"05E2", X"0589", X"0633", X"02D6", X"0011", X"022E", X"FE36", X"FE11", X"F933", X"F9F9", X"FB72", X"FCDA", X"FF9F", X"01AC", X"04B8", X"05D9", X"040B", X"0200", X"FDE7", X"FCCE", X"FC94", X"FAE6", X"FD75", X"FC38", X"FAB4", X"FA05", X"FD9D", X"02B7", X"05DA", X"0528", X"02EA", X"02CB", X"FF44", X"FFA0", X"FDE1", X"FD98", X"FCF2", X"F987", X"FA1D", X"FD9D", X"FF7F", X"025A", X"0251", X"030C", X"060E", X"05CE", X"FFE3", X"FCDB", X"FD09", X"FD2E", X"FA18", X"FC80", X"FD15", X"FF1F", X"0153", X"0488", X"04E2", X"00FA", X"02C5", X"007A", X"FE89", X"FECB", X"FD65", X"FC61", X"FB4C", X"FE76", X"FB4D", X"0007", X"FF0D", X"FE94", X"015F", X"0312", X"05F6", X"0418", X"0150", X"FEC3", X"FE35", X"FDB9", X"FE5B", X"FE6E", X"008E", X"0173", X"0161", X"031C", X"038D", X"0190", X"0109", X"FE9B", X"FDC8", X"FDC2", X"FD3B", X"FC46", X"FD29", X"FB83", X"FEAC", X"0043", X"FF6D", X"FFDA", X"00F9", X"0150", X"0200", X"0166", X"00A1", X"00F7", X"FEFE", X"FD58", X"FFBB", X"FF28", X"FFBE", X"02E2", X"FFD3", X"01C3", X"010D", X"017D", X"FE34", X"FE0B", X"FF2A", X"FE3F", X"FD3C", X"FEDE", X"FD15", X"FB51", X"FFC8", X"0079", X"FFD0", X"00A3", X"01E1", X"06B0", X"0426", X"06D2", X"041A", X"0289", X"0168", X"0206", X"011D", X"003E", X"FDB5", X"FD53", X"FF1D", X"FD9E", X"FD35", X"FEC3", X"FE6A", X"FDA9", X"FEF7", X"FC89", X"FD39", X"FF27", X"0159", X"FF12", X"FED8", X"00EE", X"0090", X"00F4", X"0161", X"068A", X"09B2", X"0895", X"0742", X"0796", X"063D", X"048B", X"042D", X"0188", X"00E8", X"FF61", X"FF45", X"FF5B", X"0018", X"0282", X"0134", X"FD8D", X"FF2B", X"01A1", X"0500", X"0446", X"FE80", X"FD78", X"FE7C", X"00F9", X"FFFD", X"005E", X"0115", X"03C6", X"0796", X"0C17", X"0697", X"0928", X"0A1B", X"0789", X"051D", X"05AF", X"0681", X"0414", X"01B8", X"00D7", X"011E", X"FF21", X"01C7", X"050A", X"0545", X"073D", X"06EB", X"0688", X"015E", X"FEEC", X"FE0B", X"00E1", X"FF24", X"FFE6", X"FFBE", X"00A2", X"0621", X"0706", X"07C8", X"07C6", X"06FF", X"0723", X"098D", X"06D6", X"08E7", X"08F2", X"08F9", X"0BBB", X"0BDD", X"09A3", X"08A9", X"0BB3", X"0791", X"05B7", X"03AD", X"00BC", X"01A8", X"00F0", X"007C", X"FFBE", X"00D7", X"003D", X"0080", X"FEFB", X"FF35", X"FF77", X"012D", X"00E7", X"0076", X"001B", X"02DC", X"02A7", X"020E", X"01AA", X"057A", X"FF9F", X"FDC7", X"01C6", X"02EA", X"FF97", X"02A0", X"0229", X"001C", X"FC68", X"0053", X"0040", X"00B7", X"0026"),
--        (X"0054", X"003A", X"FF40", X"FF8C", X"FEE4", X"FF3B", X"000A", X"0149", X"FF5C", X"FEC4", X"00E5", X"00A2", X"FDC8", X"FEE6", X"014F", X"FF91", X"FF93", X"FFE1", X"FFC6", X"00EB", X"00AF", X"FF7F", X"0038", X"FF3A", X"00EE", X"FF35", X"FF15", X"00AB", X"FFDD", X"000E", X"0067", X"00F9", X"0051", X"FE47", X"FDCA", X"FC0C", X"FD93", X"FD1E", X"FA90", X"FB0F", X"FA61", X"FB75", X"008C", X"FDF3", X"FC2B", X"FBFC", X"F957", X"FA72", X"FB1B", X"FC8F", X"FD8A", X"FD8F", X"0086", X"000F", X"FFC7", X"FF5B", X"FFEE", X"00BA", X"FE96", X"FF5D", X"FE1F", X"004E", X"FCF5", X"FC8A", X"F939", X"F881", X"F6B9", X"F740", X"F9C0", X"FC8F", X"FB89", X"FC96", X"FB09", X"FB44", X"F8BD", X"F64A", X"F6C7", X"F7DC", X"F730", X"F8F8", X"FB86", X"FD73", X"00AE", X"006B", X"FF88", X"0051", X"009F", X"FD41", X"FEB1", X"FD72", X"FB3F", X"F91F", X"F684", X"F5B8", X"F5E0", X"F6F1", X"F6BA", X"F6AD", X"F7A5", X"F7EC", X"F9EF", X"FC1F", X"FA57", X"FC02", X"F9F8", X"F932", X"F7A8", X"F624", X"F6F0", X"FB62", X"FE84", X"00BD", X"FF8C", X"FED1", X"01C6", X"FE5C", X"FFDA", X"FEC8", X"FAE5", X"F9AF", X"F81F", X"F9E9", X"F89E", X"FA64", X"FBD2", X"FB8C", X"FA66", X"F9F2", X"FD06", X"FA30", X"FD96", X"FFB9", X"FD4A", X"FCA7", X"FB03", X"FD09", X"FCFF", X"FBAE", X"FCD2", X"FBEC", X"FF01", X"00A0", X"FF3E", X"02AC", X"FF22", X"02DD", X"FDCC", X"FE70", X"FE0B", X"FC95", X"FB70", X"FB53", X"FD73", X"FC5E", X"FBF6", X"FCC8", X"FCA9", X"F9E2", X"FB12", X"FA3C", X"FB34", X"FCF8", X"FFB0", X"01D2", X"FF67", X"FBFA", X"FCCA", X"FE41", X"FFD5", X"FEE7", X"0218", X"0400", X"0222", X"0179", X"00A5", X"FF6F", X"FD44", X"FE5C", X"FE4C", X"FDD9", X"FDA8", X"FBC2", X"FE02", X"FB40", X"FB96", X"FB74", X"FB25", X"FBF6", X"FBFB", X"FBF2", X"0004", X"0275", X"02B8", X"017E", X"FECF", X"FF0E", X"0017", X"FD01", X"042D", X"0675", X"FF9F", X"FF53", X"FEDE", X"004A", X"FD7D", X"FFA1", X"FE5F", X"FE3A", X"FE97", X"FFB2", X"FD92", X"FD4F", X"FEFA", X"0175", X"0288", X"0186", X"0260", X"0264", X"025A", X"030F", X"0197", X"00ED", X"FF60", X"FE3E", X"FFDB", X"02B0", X"0491", X"025D", X"00D9", X"FE13", X"FD15", X"FEE9", X"FCBC", X"FDF7", X"FD75", X"FF23", X"FFDD", X"FEAD", X"FF89", X"02B9", X"0351", X"048A", X"04AA", X"03AA", X"0462", X"042B", X"02CC", X"01CE", X"0173", X"02AC", X"FCF0", X"FFA1", X"017A", X"03DF", X"016D", X"FF9F", X"FD65", X"FAD1", X"FB05", X"FA45", X"FC49", X"FC27", X"FE39", X"FF9E", X"001F", X"0281", X"04E9", X"0815", X"0607", X"07BB", X"0751", X"0483", X"015A", X"02CC", X"0289", X"FEDE", X"0159", X"05D7", X"0101", X"02ED", X"00B1", X"022D", X"00C1", X"0010", X"FD27", X"FAE9", X"FA94", X"FD58", X"FC64", X"FECD", X"00C1", X"008E", X"01DC", X"0189", X"03A8", X"08F7", X"060F", X"04C7", X"040F", X"03C6", X"FFB5", X"024A", X"0255", X"FFBA", X"0342", X"092E", X"078B", X"00DB", X"00AB", X"0437", X"047F", X"FD93", X"FE97", X"FD83", X"FD20", X"FEF1", X"FFB6", X"01E5", X"021C", X"0012", X"00B4", X"FEC2", X"0344", X"0839", X"04EA", X"02B8", X"01CE", X"002B", X"0113", X"020A", X"FE73", X"FCF9", X"FDEC", X"054E", X"0441", X"FF55", X"0057", X"02DD", X"045B", X"00B8", X"FF8B", X"FD07", X"00EA", X"0356", X"03A8", X"02CD", X"025A", X"018C", X"0148", X"FF10", X"021E", X"0500", X"005D", X"0199", X"FEE4", X"0010", X"FF2C", X"FD8B", X"FAB1", X"FA8F", X"F921", X"022D", X"052C", X"011F", X"019C", X"01D2", X"034A", X"01B5", X"04B2", X"0154", X"0143", X"04E4", X"03D6", X"0402", X"035F", X"FFDC", X"FDF9", X"FE45", X"020F", X"010C", X"019D", X"0227", X"FFE5", X"FFC9", X"FDF0", X"FDF0", X"FBDB", X"F6A6", X"FB6B", X"015D", X"0078", X"FE9F", X"00B4", X"0084", X"02BE", X"02B9", X"0719", X"024C", X"03F1", X"047B", X"032A", X"0486", X"FFD9", X"FC74", X"FE30", X"FDD9", X"FF96", X"00F6", X"01AC", X"0442", X"02B7", X"00E1", X"FFE3", X"FECC", X"FE26", X"FA85", X"FAEF", X"0156", X"FF89", X"FEA7", X"FFEC", X"00C7", X"016D", X"0325", X"06F3", X"02A9", X"04DC", X"04D7", X"049D", X"02CC", X"011F", X"FDC5", X"FFBE", X"FE8B", X"FF98", X"FFBF", X"03F9", X"0439", X"028F", X"FFC1", X"FECE", X"FFBB", X"FFF7", X"FE01", X"FA54", X"FEB0", X"02AF", X"00A4", X"FFA9", X"FFA2", X"FC4E", X"016B", X"03A8", X"0257", X"0575", X"06A8", X"0457", X"03B2", X"000B", X"FDB6", X"0011", X"0113", X"0100", X"017E", X"037C", X"04C5", X"01FA", X"FFDA", X"0079", X"00ED", X"FF72", X"FE6F", X"FD27", X"FB0F", X"FDFA", X"022D", X"0069", X"00D5", X"FD26", X"FE2B", X"03BE", X"049C", X"0473", X"04AA", X"04DE", X"02CB", X"01B3", X"00C7", X"0172", X"0522", X"0569", X"0526", X"016A", X"FFB5", X"FF42", X"007B", X"00D1", X"0103", X"FEE5", X"FF9B", X"FBA2", X"FF35", X"FDEC", X"FF45", X"0046", X"019B", X"FC0F", X"FF0A", X"0178", X"038F", X"0294", X"022C", X"01D0", X"022F", X"0226", X"01F7", X"02CB", X"048E", X"058D", X"0116", X"FE4F", X"FB4E", X"FDA8", X"FF53", X"FEFE", X"FD51", X"FCE5", X"FDA1", X"FAA6", X"FD20", X"00A5", X"0307", X"01AF", X"FDD2", X"FEBF", X"FE0B", X"FFD8", X"004E", X"FFE3", X"0008", X"0058", X"FF72", X"FE88", X"FFB2", X"FF35", X"FF65", X"FF68", X"FCE6", X"F95E", X"FB66", X"FC15", X"FE90", X"FCF6", X"FB58", X"FA22", X"FBDE", X"FD9F", X"0031", X"0113", X"029F", X"FF58", X"FE81", X"FC08", X"FA00", X"FAED", X"FD1A", X"FE4B", X"FD23", X"FD05", X"FAFC", X"FBAC", X"FC73", X"FA96", X"FA12", X"F9EB", X"F9C0", X"FCF5", X"FB7E", X"FAD0", X"FD33", X"FBF7", X"FC47", X"FAF2", X"FDAB", X"0131", X"02FE", X"FF8D", X"0106", X"0173", X"0172", X"FAFD", X"FAE9", X"FA2C", X"FBBA", X"F9EF", X"F86D", X"F83A", X"F89F", X"F990", X"FB4B", X"F893", X"F84A", X"FA2B", X"FA33", X"FB24", X"FAA7", X"F958", X"FBEF", X"FD3B", X"FC3D", X"FC3F", X"FCFA", X"0386", X"0525", X"FF03", X"0071", X"00B1", X"00EC", X"FCAF", X"FA5B", X"FB69", X"F8E0", X"F8B5", X"F8E8", X"FAC2", X"FB65", X"FA01", X"FC1A", X"F975", X"F967", X"FA5B", X"FA99", X"FC44", X"FBF9", X"FC71", X"FCDD", X"FD6B", X"FFE8", X"FE1F", X"0032", X"0671", X"03FF", X"030F", X"0150", X"FEF7", X"FEFA", X"FB90", X"FA15", X"FC96", X"FDB3", X"FAFE", X"FBFB", X"FC42", X"FD7B", X"FD16", X"FD2F", X"FCDC", X"FC5C", X"FDA9", X"FC63", X"FE35", X"FDEA", X"FDA1", X"0005", X"FF7F", X"FF1D", X"FF59", X"0022", X"05BB", X"04D7", X"044D", X"FFFE", X"FFBA", X"FF92", X"FDE3", X"FD78", X"001E", X"0186", X"FFEB", X"FE2F", X"FD43", X"FC7F", X"FDFF", X"FBFC", X"FBAC", X"FCDD", X"FBED", X"FBF6", X"FBE1", X"FF1F", X"FEFE", X"FF65", X"007E", X"00EA", X"0266", X"0456", X"0054", X"00A3", X"FE5E", X"0096", X"00CB", X"FF75", X"FE34", X"0427", X"0347", X"0360", X"FF09", X"FF9F", X"004B", X"FFB3", X"FCC1", X"FF23", X"FF50", X"FF5A", X"00D5", X"011B", X"FFDC", X"0031", X"019E", X"FF93", X"00DF", X"0271", X"043D", X"0531", X"044F", X"008B", X"FDC7", X"FF80", X"00E6", X"FFBF", X"00AF", X"FFED", X"FFCB", X"003A", X"01E2", X"00D1", X"0114", X"03C3", X"02D6", X"03B9", X"0285", X"03A0", X"05A6", X"0829", X"055D", X"03E5", X"04FA", X"0505", X"00ED", X"0365", X"0306", X"FFDF", X"FF67", X"00D3", X"FEF5", X"FFE3", X"FEBD", X"00C5", X"FF5C", X"FFC6", X"0046", X"FFA5", X"0138", X"FFC6", X"01CF", X"017D", X"051C", X"04E4", X"04A1", X"05A1", X"0374", X"03C3", X"0364", X"0535", X"02F4", X"0438", X"0350", X"0479", X"0353", X"0210", X"FF1C", X"006B", X"015B", X"FFBA"),
--        (X"00F8", X"008F", X"008C", X"FF2B", X"01C3", X"003D", X"002C", X"FF29", X"001D", X"006C", X"FFB2", X"FEB2", X"00E5", X"003A", X"FFBD", X"FF74", X"FF88", X"FEBA", X"0004", X"FDD5", X"FF60", X"0020", X"FF18", X"0086", X"00A3", X"0055", X"FFB2", X"0064", X"0039", X"0129", X"00D5", X"00B8", X"00AB", X"FF10", X"FF5B", X"FF62", X"FE2A", X"FDEE", X"FC79", X"02F3", X"0113", X"00F1", X"FF3B", X"0340", X"0644", X"02D1", X"FA93", X"FB76", X"FCBE", X"FE4D", X"017D", X"0082", X"FF71", X"013D", X"000B", X"FF54", X"FEFF", X"FED8", X"FFBC", X"0239", X"007D", X"FF34", X"FEB1", X"FFE9", X"FDC1", X"FEE3", X"FE87", X"FFEB", X"03B3", X"0444", X"FFAE", X"00F9", X"024C", X"FE57", X"FC7A", X"F99B", X"F8D5", X"F896", X"F857", X"FB79", X"0138", X"013D", X"FE77", X"FF7D", X"FFAB", X"FF24", X"01F2", X"0155", X"FD44", X"FC5C", X"FBDD", X"FC0A", X"FE6C", X"014C", X"FF3D", X"FF1C", X"0233", X"0306", X"0000", X"007D", X"01C4", X"FDDA", X"FAAD", X"FA08", X"F7DD", X"F524", X"F4EE", X"F52B", X"FCA4", X"FF2A", X"FD35", X"00FC", X"FF81", X"0089", X"0161", X"FF79", X"FC4A", X"FC0C", X"FF9A", X"FD56", X"FEF3", X"0047", X"FE36", X"FFA6", X"0062", X"01BC", X"04A7", X"0208", X"0155", X"FE74", X"FC1C", X"FC4C", X"FC2C", X"F76F", X"F8C4", X"F862", X"F771", X"FB79", X"01C3", X"0154", X"FFB2", X"FFD4", X"010D", X"003D", X"FD9A", X"FBED", X"FE68", X"FCA5", X"FD47", X"FD24", X"FD7A", X"FD84", X"FFAE", X"035F", X"048C", X"0565", X"0338", X"02EE", X"01EC", X"FF54", X"FFD8", X"00CA", X"FE65", X"F8A3", X"FA63", X"F917", X"FB2A", X"FC0A", X"FEE6", X"000F", X"FD7A", X"0031", X"FC62", X"FDF8", X"FE8C", X"0081", X"FD0B", X"FB49", X"FB92", X"FCE6", X"FE46", X"017B", X"01B6", X"02B1", X"02D1", X"0241", X"0195", X"0051", X"FEF8", X"011D", X"01C8", X"FDFA", X"F77F", X"F82F", X"FABC", X"FD56", X"0081", X"FB25", X"0054", X"FE76", X"0152", X"00B5", X"00E8", X"FDA0", X"FC29", X"FC3C", X"FAF1", X"FB5C", X"FD32", X"FFC5", X"014C", X"01C2", X"0403", X"0196", X"028E", X"0031", X"FEF7", X"001E", X"007F", X"FE36", X"FA57", X"F962", X"FA2E", X"FDBC", X"020C", X"FE12", X"FF5E", X"FF8E", X"031B", X"0035", X"FE90", X"FD22", X"F9B7", X"FB56", X"FCD1", X"FADB", X"FE13", X"00E4", X"0282", X"04BA", X"050B", X"043F", X"05E7", X"0347", X"00C0", X"0002", X"FFE3", X"01A6", X"FDBA", X"F92E", X"FD0B", X"FDDE", X"FFFE", X"FD50", X"0023", X"005B", X"0240", X"FE67", X"FC7A", X"F9F0", X"FA21", X"FD7D", X"FE79", X"FE93", X"FEBD", X"0192", X"025C", X"0517", X"043F", X"05E9", X"059A", X"0413", X"01C2", X"013F", X"FFF7", X"03D6", X"FF83", X"F936", X"FBC1", X"FC79", X"FFB7", X"FEB2", X"0139", X"01DD", X"FC42", X"FC09", X"FA5A", X"FB4A", X"FDA3", X"003C", X"FDF0", X"FF86", X"FCF0", X"FCA2", X"FF87", X"FF8C", X"0103", X"02D4", X"0620", X"04F3", X"04E8", X"03BC", X"04DC", X"05E5", X"047E", X"FADE", X"FDC5", X"001C", X"0026", X"00E6", X"FE04", X"FCA1", X"FB2E", X"FBDD", X"FCBF", X"FD54", X"FCF9", X"FD11", X"FBDF", X"FB5C", X"F716", X"F5DC", X"FE5E", X"FC5B", X"F994", X"FC13", X"01C1", X"044A", X"0448", X"04BD", X"045F", X"0480", X"0621", X"01F0", X"021A", X"0377", X"FF36", X"FEA0", X"FF71", X"F867", X"F9F7", X"FC11", X"FE25", X"FDDE", X"FBFF", X"FDF6", X"FAAC", X"FA4F", X"F8F3", X"FA1F", X"FE1A", X"FB35", X"F858", X"FB24", X"FE65", X"0382", X"04ED", X"0118", X"024C", X"0358", X"0659", X"05BC", X"040B", X"03BF", X"00D2", X"01C0", X"0046", X"FCA4", X"FB25", X"FC1F", X"FE9E", X"FC8E", X"FF5E", X"FF3B", X"FF50", X"FD59", X"FDF0", X"0008", X"0088", X"FBC9", X"FB39", X"FC36", X"FEDA", X"013C", X"0003", X"01E5", X"0298", X"002A", X"01E1", X"0378", X"06FA", X"0469", X"FDA2", X"FCF1", X"FECF", X"FBA8", X"FED3", X"0153", X"00C8", X"FF42", X"FF10", X"FF2A", X"FF1A", X"FF40", X"FFEF", X"03AF", X"0135", X"FD9B", X"FC1D", X"FCB5", X"FE76", X"FD48", X"00BB", X"00E1", X"FF0F", X"FF25", X"006B", X"03FB", X"08FF", X"0353", X"0004", X"FD5B", X"FDA9", X"FEE3", X"024A", X"04A5", X"00EF", X"01C9", X"01BD", X"005C", X"0145", X"FFEF", X"FE63", X"FFF9", X"FFAA", X"FFED", X"FE14", X"FBE7", X"FD7A", X"FBA6", X"FFBE", X"FF83", X"FDA0", X"FF9C", X"017A", X"04FD", X"07C1", X"03EF", X"0075", X"FB88", X"FF9F", X"018D", X"0503", X"0594", X"0481", X"0234", X"0262", X"0164", X"01CC", X"FFC5", X"FEE3", X"FFD5", X"0097", X"FFF3", X"FECC", X"FB2C", X"FCCC", X"FCD4", X"FD46", X"FF90", X"0077", X"FE47", X"0086", X"069F", X"06EC", X"031F", X"FE70", X"FCE3", X"FD57", X"04A2", X"0397", X"033E", X"037D", X"01AC", X"01FC", X"02D9", X"0468", X"00E6", X"0102", X"FEB9", X"FFA1", X"FFF7", X"FBDB", X"FA8D", X"F9CE", X"FCAE", X"FE33", X"FEF3", X"FF58", X"FDD9", X"0038", X"04CE", X"05C2", X"0301", X"0399", X"FF06", X"FA66", X"FF78", X"0195", X"0101", X"006D", X"FF73", X"00FC", X"021E", X"0287", X"0121", X"FF09", X"FF35", X"00F8", X"0023", X"FC16", X"FAF7", X"FC74", X"FB98", X"FD04", X"FF0F", X"016E", X"0084", X"02E5", X"0971", X"02E9", X"041E", X"FE3C", X"00DB", X"FA5F", X"FD31", X"0082", X"FF1E", X"FF13", X"01DA", X"00B0", X"03E0", X"0198", X"0224", X"02D8", X"0361", X"0185", X"00AD", X"FED3", X"FD09", X"FCFD", X"FD73", X"FD95", X"00C0", X"0104", X"032B", X"01E0", X"067C", X"0665", X"032A", X"FFD3", X"00AF", X"F976", X"FE4A", X"0117", X"03A1", X"0229", X"0520", X"0029", X"0123", X"0633", X"0460", X"0394", X"02A8", X"FFBF", X"008E", X"FF5A", X"FE77", X"FDD2", X"FF58", X"FF3B", X"00E1", X"032A", X"041A", X"0372", X"0372", X"02E7", X"009A", X"0023", X"FED9", X"FDC2", X"0006", X"00B5", X"02BB", X"05D9", X"03EF", X"0208", X"03D6", X"03DC", X"0108", X"FFA5", X"FF56", X"00D2", X"FF36", X"FD48", X"FD05", X"FF48", X"FE88", X"0023", X"01CE", X"0351", X"0582", X"022E", X"01C1", X"04B7", X"01C1", X"01FD", X"FECC", X"FE85", X"FE9F", X"00A9", X"04D4", X"08F6", X"0656", X"043E", X"0409", X"03A0", X"02B3", X"FFAF", X"0145", X"0073", X"FF78", X"FD60", X"FD02", X"FFC6", X"0033", X"FF4D", X"01B5", X"0281", X"01B4", X"FF3C", X"FD54", X"FD53", X"00B4", X"0054", X"FF8A", X"FCB9", X"F8BF", X"F9E4", X"FD7F", X"0029", X"01E2", X"0329", X"0415", X"0359", X"031E", X"054D", X"04AE", X"01ED", X"009A", X"0104", X"010B", X"FEC8", X"0090", X"FF29", X"011F", X"0291", X"0211", X"FD34", X"FE1F", X"FFE7", X"FFC6", X"00D8", X"FFDD", X"FDB1", X"FA21", X"F6BD", X"F786", X"F6ED", X"F90F", X"FC88", X"FCA5", X"FADE", X"FD5C", X"FF2E", X"0084", X"FEBF", X"FF08", X"FFDD", X"013E", X"0206", X"00CF", X"FE4D", X"FFFD", X"FF6B", X"FF2C", X"0477", X"0410", X"036F", X"014F", X"003E", X"FEF0", X"FFD6", X"FBE5", X"F8BB", X"F746", X"FA61", X"F879", X"F8EE", X"F648", X"F5D6", X"F7C4", X"F853", X"F8D3", X"F9A6", X"FBD7", X"FCC1", X"FC2D", X"FD77", X"FD13", X"FC06", X"FC93", X"F960", X"FC26", X"FCE1", X"01ED", X"026F", X"01C3", X"FEB3", X"FF39", X"010A", X"FE8C", X"FF6C", X"FD1A", X"FC08", X"FCBA", X"FBE4", X"F95F", X"FAFD", X"FD0E", X"FCB1", X"FC33", X"FA1D", X"F9F1", X"FA99", X"F85F", X"FADC", X"FDDE", X"FAE7", X"FA32", X"FCC2", X"FF7C", X"FF7B", X"0090", X"0093", X"FF8D", X"013E", X"FE8F", X"FF12", X"FECC", X"FEE8", X"FFB0", X"FE37", X"FFF7", X"FDE7", X"FDFA", X"FE7B", X"FE87", X"FFE8", X"FCE6", X"FED3", X"FEF5", X"FE13", X"FFD8", X"0018", X"FF52", X"FD73", X"FBE0", X"FCED", X"FE20", X"0042", X"FF95", X"FF9F", X"00FB"),
--        (X"FEA9", X"FE67", X"FF13", X"018B", X"00FE", X"0005", X"FE75", X"FFE2", X"FF81", X"0056", X"FEDA", X"0003", X"FEA7", X"FEDD", X"0033", X"0020", X"0076", X"0070", X"00D1", X"014E", X"FF65", X"005D", X"0079", X"007F", X"0168", X"FF9D", X"0068", X"FFB0", X"00CF", X"00BA", X"003A", X"FFA8", X"FEDC", X"004F", X"0061", X"FE1B", X"FF0A", X"FB61", X"F967", X"FA0F", X"FB29", X"F935", X"FFAF", X"FC45", X"FEBF", X"F95F", X"F87E", X"F9B2", X"F99D", X"FC46", X"FCA6", X"FC52", X"012E", X"0055", X"003E", X"FFB6", X"FFDD", X"FF61", X"FEB5", X"FE02", X"FBA0", X"FF37", X"FE01", X"FDB3", X"0070", X"011B", X"FF2A", X"FD08", X"F97D", X"FA29", X"FB47", X"FBBC", X"FC88", X"FBAB", X"FACE", X"F947", X"FC16", X"F893", X"F92D", X"FAAE", X"FE17", X"FFFF", X"FF94", X"0159", X"FFE8", X"FFFA", X"FF4E", X"FCFB", X"FB4E", X"020E", X"0594", X"06DA", X"07F2", X"062F", X"0404", X"04B6", X"0278", X"FFB6", X"FE40", X"FED9", X"0082", X"01FD", X"00CA", X"0013", X"00AD", X"FB5A", X"FB12", X"FA1D", X"FC21", X"FEE9", X"FF3E", X"FFED", X"0002", X"003C", X"0145", X"00BD", X"0572", X"08AF", X"0AED", X"0A01", X"0949", X"077F", X"05C1", X"042D", X"046F", X"02F0", X"FF1D", X"FCA1", X"FF10", X"FE4E", X"001C", X"FDE2", X"FCAF", X"FCCA", X"FEEC", X"FC2F", X"0142", X"FF72", X"FE2E", X"FCDA", X"0027", X"0005", X"FF13", X"0321", X"08E9", X"0CA2", X"0AB4", X"08E9", X"04C4", X"03AC", X"01FF", X"0337", X"0100", X"00A4", X"FFCE", X"FEBC", X"00E5", X"FF48", X"FF8B", X"FF31", X"FCD7", X"FE15", X"FF3F", X"001C", X"FE92", X"FF18", X"FB6E", X"FF93", X"00D3", X"00D7", X"FFF3", X"06FC", X"0A31", X"07AE", X"0869", X"03B5", X"0235", X"00C0", X"00CB", X"018E", X"FFFC", X"0087", X"FF6C", X"00D1", X"015A", X"FFE6", X"008B", X"FE9A", X"FDB6", X"FCEE", X"FDC5", X"FAE0", X"FCBE", X"FA30", X"FD10", X"FD8E", X"FF7C", X"047E", X"0172", X"070F", X"0A61", X"07A5", X"0688", X"01F1", X"0092", X"00B3", X"FF72", X"FFA9", X"004B", X"FFC9", X"00E7", X"FDCC", X"FFB9", X"FE39", X"FDE2", X"0043", X"FE7B", X"FF3D", X"FF7E", X"F980", X"F573", X"F6EB", X"FB36", X"FD07", X"FEA9", X"01D1", X"0282", X"080F", X"0AEB", X"084D", X"0577", X"02F4", X"0088", X"FCE9", X"016C", X"FDB8", X"FDFC", X"FFC5", X"FE89", X"007A", X"017C", X"0186", X"FFDA", X"FFC8", X"0156", X"FFFD", X"FE4D", X"F900", X"F228", X"F5DF", X"F953", X"FDD7", X"00EC", X"02F5", X"0237", X"05A1", X"0AA7", X"0869", X"06A1", X"0352", X"FE14", X"FD38", X"FDDE", X"FAAD", X"FC21", X"FD07", X"0078", X"0572", X"0765", X"06E4", X"0460", X"0368", X"02E7", X"005B", X"026F", X"F9F4", X"EF30", X"F3CC", X"F779", X"FD5B", X"FF7C", X"0203", X"00D4", X"0819", X"06F9", X"08D8", X"03E1", X"FEDD", X"FB81", X"F82A", X"FAB1", X"F953", X"FC37", X"FB8F", X"FD10", X"038C", X"0608", X"0657", X"04C4", X"0583", X"02AC", X"023A", X"034D", X"F9FE", X"ED1D", X"F5EC", X"FD28", X"FEAC", X"FFB1", X"00B7", X"0382", X"0776", X"0913", X"0546", X"FEBD", X"FB0E", X"FAF1", X"FB42", X"FD92", X"FDDC", X"FDDB", X"FA68", X"FC5F", X"02A5", X"0579", X"05FA", X"03B8", X"05C1", X"0305", X"FFAB", X"009B", X"F9E1", X"EE37", X"F6E3", X"FD9C", X"FF7C", X"FFCD", X"02B0", X"03BF", X"0240", X"056D", X"0302", X"FD67", X"F928", X"FE5D", X"FDE2", X"0142", X"0065", X"FEDC", X"FABE", X"FBC2", X"FFCE", X"047F", X"02DF", X"040D", X"03EF", X"FF88", X"FDA5", X"FC55", X"F633", X"F6CB", X"0228", X"060B", X"0334", X"FF1C", X"FF29", X"0336", X"00A9", X"03D7", X"00EE", X"FDD6", X"FD71", X"0014", X"00C6", X"026D", X"FF0D", X"FD19", X"FE4B", X"FE9C", X"0032", X"0455", X"0406", X"03A5", X"0283", X"00F0", X"FE2C", X"F932", X"F806", X"FB73", X"03BE", X"08FC", X"0426", X"FDE4", X"01F4", X"0039", X"03D1", X"0220", X"00D7", X"005A", X"0090", X"004D", X"FF7B", X"FE68", X"FCE6", X"FD87", X"FC4B", X"FE4B", X"0114", X"0472", X"03B0", X"047A", X"046F", X"0108", X"FFD3", X"FE90", X"FA6F", X"FC95", X"023A", X"0840", X"029C", X"FD45", X"0045", X"024B", X"0692", X"03DF", X"0311", X"0401", X"00C5", X"FF2A", X"FD98", X"FA0A", X"FDC1", X"FCA5", X"FC5E", X"018B", X"05C3", X"05B5", X"04D0", X"01E5", X"04D6", X"02F1", X"0265", X"02F2", X"FF3A", X"014B", X"0488", X"0B19", X"02B9", X"0184", X"0179", X"02A2", X"04E6", X"06A6", X"0573", X"0369", X"00C4", X"FC9A", X"FC4C", X"FC6A", X"FC9F", X"FD3D", X"FFB1", X"0482", X"0599", X"0676", X"04ED", X"044F", X"04F0", X"0192", X"02AB", X"0255", X"012E", X"030A", X"0651", X"0C17", X"038C", X"FFE5", X"01BB", X"03C6", X"06C8", X"05FE", X"026B", X"0218", X"019F", X"FE01", X"FAA0", X"FA8F", X"FC56", X"FEA7", X"0136", X"0614", X"07F7", X"06B5", X"0333", X"052E", X"026C", X"0134", X"0176", X"0132", X"02A8", X"0332", X"07C8", X"09AF", X"0115", X"00F2", X"0187", X"0259", X"05BC", X"06BA", X"03EF", X"024C", X"FEEE", X"FCD4", X"FA09", X"FB7C", X"F928", X"FCBE", X"0429", X"06F4", X"0413", X"0545", X"037A", X"063C", X"03A5", X"00F9", X"01A4", X"020A", X"02C4", X"002E", X"070E", X"0713", X"03AA", X"0051", X"FED0", X"FEDD", X"0337", X"0432", X"02A9", X"014A", X"FE29", X"FD0F", X"FB81", X"FA60", X"FA90", X"FC0F", X"013C", X"030F", X"0387", X"03E0", X"02A8", X"027E", X"0185", X"00CF", X"0140", X"FD5F", X"01CD", X"023D", X"054F", X"04CD", X"00EF", X"FF3D", X"FE70", X"FD97", X"02CF", X"03DA", X"014F", X"014D", X"FEFC", X"FCEF", X"FB9F", X"FA2C", X"F86C", X"FA0C", X"FCDE", X"FF9C", X"FE9D", X"010B", X"0181", X"01D8", X"010C", X"0099", X"FDF9", X"FE0E", X"FFD6", X"02EF", X"056A", X"05C2", X"FE7A", X"FD64", X"0252", X"049C", X"01EA", X"00B0", X"FE0E", X"FE73", X"FCD8", X"FD8D", X"FC2F", X"FC9C", X"FB13", X"FBC7", X"FBBA", X"FBB0", X"FDCA", X"0076", X"FFB8", X"0092", X"0161", X"FE6A", X"FD4F", X"01A1", X"0235", X"020E", X"0111", X"00F2", X"FF6A", X"0033", X"FF70", X"0734", X"02D1", X"00A2", X"FE36", X"FFD9", X"FCFF", X"FE5E", X"FE1E", X"000F", X"FE0D", X"FEFB", X"FD7F", X"FBB7", X"FDAC", X"FE3E", X"FF4E", X"007F", X"FF6E", X"0360", X"0172", X"04A1", X"031B", X"02DF", X"0055", X"FDF6", X"FFE5", X"FFB8", X"00A0", X"FFFD", X"0439", X"0167", X"FE9A", X"FF0B", X"FF5C", X"FC0A", X"FCD4", X"FF2C", X"FFAF", X"FE5C", X"FEA4", X"FE37", X"FF1F", X"FD9C", X"FEA2", X"0149", X"00D9", X"0550", X"0604", X"057D", X"FF59", X"013D", X"0027", X"0159", X"FF6A", X"0105", X"FFD0", X"024F", X"03C5", X"0616", X"039B", X"03AE", X"03A8", X"0057", X"FF3E", X"FF0D", X"FFD0", X"FDF9", X"0007", X"003A", X"FF03", X"FFB5", X"00F0", X"0064", X"0093", X"0327", X"04CA", X"036A", X"FF4D", X"FF30", X"037D", X"04D0", X"007F", X"00B3", X"0063", X"00D6", X"FE91", X"05CA", X"0964", X"0901", X"0712", X"07E9", X"03B0", X"028A", X"FF37", X"0262", X"0056", X"00FD", X"00AC", X"016C", X"FFCA", X"FF3F", X"0041", X"01FA", X"FF79", X"FCDC", X"FBD6", X"FC75", X"01B1", X"0328", X"0075", X"0058", X"FFEA", X"0008", X"0186", X"01B0", X"0293", X"05D0", X"05DB", X"063A", X"04E9", X"048C", X"0062", X"0024", X"0265", X"0584", X"068A", X"03A6", X"044C", X"0297", X"01E8", X"003F", X"FED0", X"FF96", X"0089", X"FF6E", X"FF8B", X"FF55", X"0062", X"FF21", X"0009", X"FF9B", X"FFCC", X"FF69", X"014A", X"014F", X"0235", X"0101", X"01B1", X"00A9", X"FED6", X"FF82", X"034A", X"04F1", X"0259", X"013E", X"021C", X"01DB", X"0252", X"0355", X"02A3", X"0304", X"00C6", X"FE9B", X"FEF2", X"FFA7", X"FEDB"),
--        (X"009D", X"FEFB", X"FFD7", X"010C", X"00B5", X"FF76", X"0044", X"FF7B", X"FFEB", X"00CD", X"0026", X"FFBD", X"FFEF", X"0085", X"FFD6", X"0014", X"FEC2", X"FF7F", X"0026", X"0087", X"FE77", X"FFF9", X"FF6D", X"FF75", X"FF43", X"008D", X"FFE4", X"FEA5", X"FFC6", X"FF17", X"0108", X"0016", X"003B", X"FFFC", X"FD33", X"FBAE", X"FCC5", X"FDAD", X"FD13", X"FBD7", X"FABE", X"FC58", X"FFB3", X"FCDA", X"FBAB", X"FC7B", X"FC4B", X"FC95", X"FC52", X"FCA7", X"FD23", X"00C6", X"FE8F", X"FE59", X"004E", X"00B9", X"008E", X"00D5", X"FF51", X"FCB5", X"FE5E", X"FEED", X"FC56", X"FB58", X"F996", X"FA86", X"F7C5", X"F695", X"F8CE", X"FCA2", X"FB59", X"FA12", X"F97D", X"FB48", X"FB38", X"FCB7", X"FC67", X"FB1D", X"FC29", X"FAED", X"FB34", X"FC4A", X"0102", X"00C5", X"016E", X"00B2", X"01E0", X"FD83", X"FE0B", X"FAAD", X"FB03", X"F9A7", X"F7EE", X"F894", X"F9E3", X"F6CD", X"FB37", X"FB28", X"FB50", X"FCF8", X"FA42", X"FA42", X"FC51", X"FE58", X"FE14", X"FF43", X"01F6", X"FF42", X"FBE9", X"FF05", X"0075", X"00C9", X"FE8D", X"FEDC", X"01CD", X"FC6D", X"00AA", X"FBB0", X"FBD4", X"FDE0", X"FD4D", X"FBB1", X"FB1A", X"FE98", X"FEC8", X"FE80", X"0085", X"FF88", X"FECC", X"0071", X"0010", X"FFEE", X"0154", X"030D", X"039B", X"044E", X"0538", X"0278", X"0111", X"FDCD", X"002C", X"020E", X"00B0", X"FCAB", X"FC5F", X"FC85", X"FD67", X"FE7C", X"FBF0", X"FE96", X"FE89", X"FFB2", X"0183", X"FF69", X"FF30", X"FF7E", X"FE37", X"FE04", X"FEF6", X"FF17", X"0171", X"0238", X"0341", X"04E4", X"0233", X"0348", X"0362", X"FDE3", X"0009", X"FE3C", X"FEF9", X"FB33", X"FCF0", X"FC0D", X"FDF8", X"FEE9", X"FE7B", X"FF01", X"FE72", X"FF7C", X"FF27", X"FD15", X"FF5A", X"FF3D", X"FDB3", X"FF24", X"000F", X"01B6", X"01B5", X"00B8", X"01B4", X"06FC", X"06B3", X"0716", X"08C5", X"0449", X"FF97", X"FD94", X"FE14", X"FA40", X"F97E", X"FB66", X"FBD2", X"FD6F", X"FD88", X"FB7D", X"FDF5", X"FDAD", X"FEBC", X"FE3B", X"FD36", X"FCFC", X"FFD8", X"FCED", X"00FD", X"0109", X"0261", X"0162", X"02D2", X"0500", X"0578", X"0553", X"0966", X"028F", X"FE31", X"FD3D", X"FEDA", X"F9AB", X"F7D9", X"FA53", X"FBEB", X"FD9F", X"FE80", X"FF05", X"005A", X"026D", X"0318", X"007A", X"FC80", X"F98B", X"FBAB", X"FDFF", X"FCFC", X"FE59", X"FFFF", X"0021", X"00FF", X"045D", X"09FD", X"0A4F", X"0A1D", X"03EF", X"FFBF", X"0088", X"FE70", X"FB4F", X"F9C4", X"FC19", X"FE97", X"01FF", X"0387", X"0292", X"04F7", X"07B9", X"0639", X"016A", X"FCA4", X"F983", X"F7BF", X"FB6D", X"FBED", X"FCB0", X"FD89", X"FF07", X"003C", X"FFC8", X"07DF", X"0733", X"08D1", X"027E", X"FEEE", X"FFC6", X"FE6C", X"FC0C", X"017E", X"02CE", X"056F", X"0930", X"093A", X"09DF", X"0AF0", X"0A47", X"09F3", X"055D", X"FFCD", X"FFD5", X"FD3C", X"FB98", X"FC9A", X"FCC6", X"FA63", X"FD88", X"FBE9", X"FC2B", X"035B", X"0864", X"0795", X"029F", X"FF4E", X"FD0F", X"FF6B", X"FE74", X"0502", X"0A09", X"0BBC", X"0E25", X"0AC3", X"0A1F", X"0856", X"0721", X"04FC", X"039D", X"05B3", X"034A", X"01F8", X"0129", X"FF97", X"FDE0", X"FB9C", X"FC91", X"FD55", X"FDFD", X"025C", X"070D", X"083B", X"024B", X"FF8B", X"00DC", X"016F", X"04A7", X"0BCD", X"0D47", X"0D9A", X"0CFD", X"0820", X"055A", X"041D", X"0268", X"0019", X"00E6", X"04AA", X"079B", X"03E5", X"0252", X"00F2", X"00E0", X"01A6", X"FFDB", X"FD68", X"FB2E", X"FE33", X"0033", X"00C6", X"009E", X"0001", X"0145", X"00FB", X"04B0", X"09FC", X"0817", X"0728", X"03CA", X"003D", X"0039", X"000B", X"FE70", X"FD52", X"01E6", X"0430", X"0627", X"0656", X"0271", X"0143", X"054D", X"035D", X"0094", X"FD89", X"F992", X"F882", X"FAE4", X"FD05", X"FD67", X"00CE", X"00DC", X"0091", X"0323", X"045D", X"01B0", X"FF2F", X"FD75", X"FE06", X"FD54", X"FEBC", X"FD5F", X"FE4E", X"00B8", X"03D6", X"052F", X"0398", X"02D4", X"0363", X"0551", X"01D0", X"FF59", X"FD72", X"F9BC", X"F621", X"F9BD", X"FAB2", X"FDE7", X"0120", X"FE3D", X"FE4C", X"02B4", X"FF46", X"FA40", X"FBE6", X"FA20", X"FB7E", X"FCD5", X"FF21", X"0069", X"0053", X"013A", X"02ED", X"02D4", X"021A", X"0091", X"0243", X"0241", X"FFC6", X"FF08", X"FCF5", X"FAC9", X"F52C", X"F53C", X"F737", X"FD0B", X"FF81", X"FE54", X"FCAB", X"FDF4", X"FBB6", X"FAD2", X"FAA9", X"FB4A", X"FE16", X"FD61", X"FF8E", X"FF5A", X"0076", X"00B8", X"0448", X"02F7", X"003A", X"FF94", X"FF2B", X"FF66", X"FE48", X"FEC7", X"FEF9", X"FB9B", X"F6AB", X"F3A1", X"F8BD", X"FCE4", X"FF80", X"FFF2", X"FBE7", X"FA91", X"FB79", X"FC4F", X"FC23", X"FC41", X"FD8E", X"0058", X"01A4", X"03BB", X"01BD", X"0435", X"03B4", X"032F", X"FF62", X"FE68", X"FFA1", X"FD16", X"00D1", X"FF5A", X"FDEE", X"FFA1", X"FDE4", X"F720", X"FBAB", X"FC3E", X"FED9", X"FED5", X"FD69", X"FAA5", X"F9B6", X"FD04", X"FE25", X"FEE9", X"FD4D", X"FFCD", X"0194", X"028F", X"0355", X"057A", X"05D8", X"01DD", X"FCF5", X"FC3E", X"FC51", X"FFB0", X"00FA", X"FFE9", X"FEA3", X"FFA9", X"00B8", X"F900", X"00B1", X"FD06", X"01D8", X"FD4D", X"FDEB", X"FB91", X"F988", X"FE45", X"FFA4", X"FD22", X"FD45", X"FEEB", X"FE0F", X"FD4B", X"00CC", X"010A", X"0148", X"FDD7", X"FC84", X"FC4A", X"FD87", X"FEAB", X"010D", X"FEE7", X"FF06", X"00B6", X"01FE", X"FB5E", X"FF87", X"008F", X"FF8B", X"FDF4", X"FB45", X"F8CD", X"F9C3", X"FE4B", X"FCF1", X"FB97", X"FE00", X"FB9A", X"FE38", X"FD6E", X"FEFE", X"FDD8", X"FDD1", X"FD5B", X"FF15", X"FF25", X"002E", X"FF82", X"FEB6", X"FFDC", X"01F0", X"0575", X"0040", X"FD7C", X"007E", X"0138", X"01E2", X"FE9A", X"FA2F", X"FAA1", X"FCAB", X"FFE8", X"FF8C", X"FD5A", X"FEDF", X"FF7F", X"FE60", X"FE89", X"FDB3", X"FD01", X"FEDE", X"FF6F", X"FFAC", X"FF96", X"FE8D", X"FF32", X"026C", X"033E", X"042F", X"008A", X"FEE9", X"FE30", X"FB9F", X"006E", X"0062", X"FF79", X"FB93", X"FAFD", X"FE86", X"FF77", X"FEB5", X"FFFC", X"FE88", X"0020", X"FE5F", X"FEEE", X"FF34", X"0026", X"FECE", X"FDAE", X"FE26", X"FF30", X"FF83", X"FE5F", X"FF98", X"013C", X"0154", X"0181", X"00F7", X"018E", X"0133", X"FF0B", X"000C", X"FF2F", X"FC68", X"FACF", X"FD3B", X"0053", X"FD33", X"FE6F", X"FEA5", X"FE20", X"FE82", X"FE2B", X"FFB1", X"00BD", X"FE77", X"FF30", X"FF69", X"FDD8", X"FE2F", X"FF6B", X"0163", X"0133", X"FEB5", X"017F", X"00DA", X"0168", X"01B9", X"FE99", X"00DC", X"001F", X"FD52", X"FAC2", X"FA82", X"FF15", X"FE17", X"FE29", X"FFDA", X"0069", X"FF54", X"FF23", X"FFA1", X"FC57", X"FDC8", X"FFF0", X"FD28", X"FE9C", X"020D", X"03A8", X"0226", X"FFFE", X"FECE", X"02CC", X"FD23", X"FE55", X"FF7B", X"0016", X"FFAA", X"FF5A", X"FFB8", X"0355", X"FF85", X"FF2C", X"FDCF", X"FF73", X"FE36", X"FE2F", X"FD8E", X"FD03", X"FD06", X"FCE2", X"FF08", X"FFE8", X"FEB8", X"FDBA", X"003D", X"007C", X"02E4", X"03AE", X"00CA", X"04B7", X"0402", X"FE30", X"FF20", X"0116", X"0089", X"FF8A", X"FF95", X"001E", X"0107", X"04DC", X"0533", X"0139", X"017B", X"06AA", X"011D", X"00B7", X"0031", X"015A", X"01B8", X"0116", X"FEE0", X"FF06", X"FEDA", X"FEBA", X"0185", X"003A", X"FFF9", X"007B", X"00C3", X"FF21", X"0064", X"FFB6", X"FF58", X"00BB", X"003F", X"010E", X"FFCC", X"00A8", X"0193", X"020F", X"021B", X"0185", X"0315", X"031D", X"0479", X"031C", X"0346", X"01FF", X"0221", X"01DE", X"02EF", X"0278", X"0085", X"00A7", X"01FB", X"FF8B", X"FF77", X"FFF8", X"FE79", X"0002"),
--        (X"0035", X"FFE5", X"FEAB", X"002E", X"FEFC", X"0063", X"FF61", X"0026", X"00A3", X"000D", X"FFBA", X"009E", X"0052", X"FEBD", X"FF91", X"FFEC", X"FFA5", X"FF3E", X"FF2A", X"FE87", X"00C2", X"003D", X"005C", X"FFE7", X"0199", X"0010", X"FEB7", X"003E", X"005C", X"FF1D", X"0079", X"FF5E", X"FFA0", X"0165", X"03B4", X"0388", X"0499", X"040E", X"0668", X"0343", X"0360", X"037A", X"0156", X"024D", X"0363", X"04F5", X"052E", X"068E", X"06B7", X"042A", X"0407", X"011E", X"0084", X"FF1D", X"0100", X"004D", X"01FF", X"0054", X"008F", X"009F", X"017A", X"0349", X"044E", X"082A", X"0840", X"0B11", X"0A9E", X"0B66", X"0BC9", X"0A21", X"09F7", X"0A08", X"07F5", X"0853", X"09E4", X"098E", X"0947", X"085A", X"07AD", X"0620", X"0211", X"013B", X"FEA0", X"FE81", X"005B", X"00C8", X"002D", X"031F", X"0603", X"032F", X"05C9", X"075C", X"0852", X"0BA8", X"0A5D", X"0CCF", X"0E61", X"0C6A", X"0798", X"058A", X"04FC", X"060B", X"065B", X"07BA", X"06B8", X"052C", X"02CB", X"0285", X"029F", X"FF6A", X"02DC", X"0111", X"0081", X"0096", X"FFD5", X"00D7", X"0376", X"041F", X"02D4", X"02F4", X"0664", X"0756", X"06EA", X"064C", X"048D", X"027B", X"FDF3", X"FEC6", X"FFF1", X"FFD0", X"01C1", X"012E", X"00FC", X"02C1", X"0269", X"0317", X"023E", X"FF21", X"FE94", X"FFE2", X"FF27", X"FFEB", X"03BD", X"020D", X"059C", X"0128", X"01A0", X"0242", X"0442", X"02F8", X"043B", X"00BE", X"FE1F", X"FF4F", X"FDCD", X"0045", X"FFC4", X"FBD9", X"FEA9", X"0015", X"FFD0", X"012B", X"01A5", X"0479", X"040B", X"00E9", X"039E", X"02EF", X"0142", X"FFC6", X"0306", X"0194", X"0551", X"0003", X"FEF1", X"00A3", X"012D", X"0147", X"0124", X"005E", X"006A", X"FF19", X"FF5C", X"FEBC", X"FCB0", X"FDED", X"FE63", X"FD4C", X"FD93", X"FCBF", X"FD41", X"004D", X"0571", X"04F2", X"050A", X"0184", X"000E", X"01E9", X"0188", X"FF0A", X"042D", X"00E4", X"FF12", X"FEFF", X"FDF5", X"FD93", X"FF3B", X"FDBA", X"FE95", X"FD5B", X"FED9", X"FC11", X"FAFF", X"FB4E", X"FAF1", X"FD22", X"FB2C", X"FC7C", X"FD66", X"FEE3", X"039D", X"0824", X"057F", X"FFB8", X"FD80", X"009C", X"FF49", X"FEE2", X"021F", X"FF43", X"F8F1", X"FBD8", X"FD8F", X"FCFF", X"FDD2", X"FB9A", X"FB19", X"FA6D", X"FEA8", X"FC8F", X"FD03", X"FC2C", X"FB20", X"FB00", X"FCEA", X"FC6A", X"FE21", X"FF96", X"0500", X"0798", X"02DF", X"FF27", X"FED7", X"FDDA", X"FD39", X"FE3D", X"0087", X"FBA5", X"F98F", X"FC1A", X"FE55", X"FB2C", X"FA79", X"FAA8", X"F98E", X"FAC6", X"FC85", X"001C", X"FF37", X"FD64", X"FB35", X"F881", X"FC20", X"FEB0", X"FE7E", X"FE68", X"048F", X"08C7", X"0481", X"01AD", X"0054", X"01E8", X"FDEE", X"FDC5", X"FCEA", X"FB6E", X"FA99", X"F9FC", X"FB55", X"FAFE", X"FB13", X"FA89", X"FB34", X"FF78", X"FFA8", X"0249", X"0235", X"FE21", X"FC2F", X"FA91", X"FDC6", X"FDDD", X"FD07", X"0127", X"06D6", X"0BF2", X"04CF", X"0117", X"FFEC", X"FDB3", X"FF17", X"0048", X"FC43", X"FB9B", X"FABA", X"FC9F", X"FAC1", X"FA0F", X"FC7B", X"FD36", X"FE8E", X"01BA", X"02F8", X"0339", X"0186", X"0055", X"FE67", X"FD8A", X"FD75", X"FC03", X"FB02", X"F968", X"FF61", X"0724", X"01BD", X"00F1", X"002D", X"FCFA", X"FBAD", X"FF78", X"FDAC", X"FEAB", X"FDC7", X"FDD0", X"FE1F", X"FD15", X"012F", X"02DE", X"0442", X"0324", X"0264", X"034F", X"005A", X"005A", X"FDE7", X"FCE9", X"FD3F", X"FB5A", X"F7B9", X"F876", X"F8B7", X"FFD8", X"03F0", X"FF69", X"FFD7", X"FE9C", X"FCA1", X"01CC", X"FED9", X"FFEE", X"FFA1", X"FE9A", X"0161", X"0207", X"0317", X"0130", X"0237", X"04C0", X"02D9", X"01CA", X"FFBE", X"FE3F", X"FE05", X"FD42", X"FDEA", X"FCBE", X"FD81", X"FDCF", X"FEE8", X"014E", X"0041", X"FD31", X"01BA", X"01B2", X"FFA7", X"041C", X"FFC3", X"FEA4", X"FF9D", X"FFF2", X"FF9C", X"01CC", X"0157", X"0056", X"0315", X"02B6", X"025E", X"00A9", X"010D", X"FEF3", X"0040", X"0164", X"FEF2", X"00D0", X"01E0", X"01D3", X"02BA", X"011E", X"00E6", X"FECE", X"021E", X"0144", X"0462", X"0458", X"FF38", X"FD59", X"FCDC", X"FC58", X"FADE", X"FC0B", X"FD79", X"FF8F", X"FFEB", X"0178", X"015F", X"FDA9", X"FCC7", X"FDCC", X"0209", X"023F", X"01AD", X"010D", X"03AA", X"04D4", X"0728", X"03A5", X"FA70", X"FF34", X"0025", X"0220", X"042B", X"07FB", X"02EC", X"FF12", X"FD7A", X"F9B1", X"F753", X"F7CC", X"FAA1", X"FC7D", X"FEBF", X"0169", X"0112", X"FD03", X"FCE2", X"FDA2", X"0279", X"04DF", X"02E6", X"01A4", X"032C", X"043E", X"0602", X"0372", X"FEC7", X"FDC9", X"0022", X"0330", X"0201", X"083C", X"0392", X"027E", X"FF53", X"FA6A", X"F9C2", X"F88F", X"FC6B", X"FA94", X"FBA2", X"FFB4", X"FF0E", X"FBAC", X"FE1F", X"FEA8", X"0126", X"0404", X"02F0", X"03A7", X"02BC", X"0474", X"0242", X"03FC", X"0035", X"FCFF", X"FECC", X"00CA", X"048F", X"08FE", X"0366", X"0142", X"024A", X"00BA", X"FFB6", X"FF4F", X"FF31", X"FE3D", X"0286", X"0385", X"01C6", X"FEA9", X"006F", X"0204", X"0194", X"03EB", X"048F", X"048B", X"03BE", X"0444", X"02B3", X"0841", X"00EE", X"02BA", X"0080", X"FE5C", X"0331", X"0583", X"0315", X"012E", X"02BA", X"037D", X"0485", X"054A", X"02CA", X"0555", X"0462", X"05A8", X"0447", X"02C0", X"04DF", X"04A4", X"0391", X"0398", X"02EB", X"052B", X"0157", X"021B", X"024E", X"0492", X"FFA8", X"02C1", X"FFC1", X"FE00", X"0180", X"0637", X"0076", X"FFB5", X"029F", X"04EF", X"05CC", X"0690", X"0724", X"068A", X"04AE", X"03B3", X"043A", X"030A", X"0448", X"01E2", X"0440", X"02D6", X"02B1", X"0121", X"015B", X"FFCF", X"0299", X"04CE", X"0262", X"0062", X"01AB", X"010F", X"0335", X"0359", X"00A6", X"0140", X"041C", X"0523", X"0388", X"0409", X"0547", X"017A", X"0088", X"FF6B", X"0204", X"02F0", X"01C6", X"0241", X"03D8", X"0172", X"01B6", X"0152", X"FFBD", X"FF25", X"03DB", X"053D", X"024A", X"0018", X"018C", X"FF69", X"0361", X"01D7", X"01E7", X"01B9", X"0129", X"0032", X"0001", X"0371", X"0095", X"FE6F", X"FE24", X"FD6E", X"FD99", X"FF5A", X"0177", X"FF36", X"006B", X"000C", X"FF9D", X"0050", X"FC52", X"FE85", X"FFA7", X"039D", X"0277", X"0052", X"00B3", X"01F6", X"027B", X"0487", X"062A", X"05B8", X"02DB", X"FFED", X"FFC3", X"0175", X"00F8", X"FE66", X"FD0D", X"FBB9", X"FB71", X"FBC2", X"FC46", X"FD46", X"FD5F", X"FDE7", X"FEA8", X"FCD3", X"FD80", X"FDC3", X"FFBA", X"034B", X"04C0", X"FE87", X"00CE", X"0089", X"FFCE", X"03E4", X"025F", X"0262", X"0115", X"FFE5", X"FF53", X"00E9", X"0170", X"FDBE", X"0037", X"FE65", X"FD7E", X"FBD0", X"F8D5", X"FC9C", X"FA23", X"FA5B", X"FBA5", X"FDBF", X"FEA6", X"FC55", X"FFEE", X"045F", X"025B", X"FED4", X"0072", X"FEB0", X"0142", X"FF12", X"FD92", X"FC65", X"FDBF", X"FCE5", X"FCBB", X"FD00", X"F93D", X"FA9A", X"FD59", X"FBF9", X"FAD2", X"FAE7", X"FB07", X"F99A", X"FA15", X"FEA0", X"FCFE", X"0008", X"0071", X"FF8D", X"FFCB", X"00A7", X"FFDA", X"FFC4", X"000A", X"0111", X"FF8D", X"0145", X"FE37", X"FCB0", X"FC42", X"FB32", X"F935", X"FA5F", X"F8E9", X"F8EB", X"F977", X"FA2B", X"F962", X"F9D8", X"F9B9", X"FB35", X"FD8E", X"005E", X"023B", X"0274", X"0260", X"FE7E", X"FFE2", X"00AC", X"FF5F", X"FFAA", X"0112", X"FFBA", X"00F6", X"0055", X"0016", X"FF40", X"FF74", X"FE28", X"FF07", X"FDF6", X"FCB1", X"FD19", X"FDAA", X"FDEA", X"FF0B", X"FE24", X"FE2B", X"FDF3", X"FF3B", X"FD8D", X"FF57", X"FD75", X"FF4D", X"0113", X"FFD6", X"0125", X"FE42", X"FF89"),
--        (X"0102", X"FF89", X"004B", X"FFA5", X"0025", X"FF6F", X"FF72", X"0103", X"FF34", X"0021", X"FF4E", X"008B", X"FF75", X"FE8E", X"FF41", X"0119", X"FF77", X"FF1A", X"0039", X"007A", X"FFAE", X"00CA", X"00D9", X"00C2", X"FF45", X"FFF0", X"FF4E", X"00E0", X"FF7F", X"FF19", X"0006", X"FF67", X"0008", X"FEAC", X"FBEB", X"FC3F", X"FB6B", X"FDFD", X"FC86", X"FBC9", X"FB45", X"FBDB", X"FEAB", X"FBD4", X"FC55", X"FCB1", X"FE28", X"FD5D", X"FCC2", X"FDF7", X"FCFF", X"FD9A", X"FF90", X"0049", X"0067", X"00C5", X"00CC", X"006C", X"FE9E", X"FF16", X"FDD7", X"FF21", X"F9DA", X"FAF3", X"F987", X"F85A", X"F904", X"F929", X"F971", X"F7E3", X"FA0A", X"FBD4", X"FB8B", X"FC6A", X"FD7E", X"FE7E", X"FCE4", X"FCA0", X"FBB1", X"FC03", X"000C", X"FF93", X"FFF2", X"FF59", X"00B3", X"FF10", X"0194", X"FDAF", X"FE2E", X"00B9", X"FCEE", X"F898", X"FA6E", X"F8A5", X"F782", X"F969", X"F733", X"F528", X"F774", X"F89D", X"F9E4", X"FBF5", X"FEBD", X"FF04", X"FAB6", X"FA74", X"FE4B", X"FDA7", X"006A", X"FFA7", X"FFE4", X"FF18", X"014A", X"0143", X"00AC", X"0360", X"0116", X"FEC2", X"FD9E", X"FD9A", X"FDAA", X"F90F", X"FA1F", X"FAAA", X"F92F", X"F9B4", X"F964", X"F891", X"F8B1", X"F8C7", X"FC86", X"FA8A", X"FA04", X"FCA4", X"FBCB", X"FB7E", X"0074", X"FFFD", X"FE50", X"FF43", X"FF63", X"FF88", X"FF65", X"02CA", X"02C2", X"0239", X"0008", X"01E4", X"00FC", X"00A5", X"FDEA", X"FFC0", X"FEB7", X"FC57", X"FC7B", X"FEA9", X"FD22", X"FD54", X"FCAD", X"FB12", X"FBBD", X"F9ED", X"F98A", X"FA63", X"FD8D", X"FE3C", X"FAE2", X"FED4", X"002E", X"FFC3", X"0164", X"03DE", X"01D1", X"028D", X"0042", X"008F", X"024A", X"0314", X"04AE", X"01C5", X"0164", X"0294", X"01C3", X"0080", X"01C4", X"0204", X"0135", X"FE12", X"0062", X"0007", X"FE0E", X"FAD0", X"F9A7", X"FBD3", X"FD51", X"FF5B", X"FF13", X"0448", X"0242", X"03B1", X"01C5", X"00B8", X"012D", X"009D", X"0280", X"0237", X"02E9", X"02D6", X"0413", X"039D", X"028D", X"0311", X"0413", X"04C2", X"021B", X"FF75", X"01BD", X"FF3F", X"FCF4", X"FE43", X"FEB9", X"FD52", X"FF1D", X"0089", X"FCD8", X"01FF", X"0218", X"04B9", X"01B4", X"FF11", X"0025", X"01AB", X"0265", X"00F4", X"0055", X"00C4", X"0227", X"FFA6", X"0147", X"0129", X"00FF", X"00F6", X"0033", X"FF51", X"FF3B", X"FFE1", X"004E", X"FFFF", X"FEC5", X"FEED", X"FD43", X"FD7D", X"00AC", X"02FC", X"008B", X"02B2", X"00CA", X"00FC", X"00FE", X"0072", X"041D", X"0119", X"001B", X"FFDE", X"0206", X"032F", X"0242", X"01D6", X"015B", X"FE4A", X"001D", X"FFF3", X"0052", X"0128", X"0093", X"FDE5", X"FE52", X"FECF", X"FB37", X"01DA", X"01E0", X"013A", X"024F", X"04E4", X"010A", X"FF91", X"FFC4", X"FFB2", X"FF44", X"FF38", X"0051", X"0231", X"0293", X"FF9C", X"FE7C", X"028A", X"0298", X"FF78", X"FF60", X"FFC4", X"0048", X"0146", X"0035", X"FD00", X"FCDA", X"009C", X"FBD2", X"0094", X"00DA", X"0098", X"0527", X"0823", X"0311", X"FECE", X"FE8B", X"FE8B", X"FED0", X"0015", X"02BB", X"0475", X"FEC7", X"FB3D", X"FE1F", X"025F", X"031C", X"02CC", X"01A1", X"000B", X"030B", X"006D", X"0146", X"FB3D", X"F898", X"0009", X"FCA1", X"FFC7", X"0054", X"0243", X"0478", X"03D5", X"020F", X"0096", X"FF2B", X"FE1A", X"FED7", X"FEAD", X"03DB", X"0217", X"FC94", X"FCF4", X"01BB", X"04B2", X"0461", X"029D", X"02D5", X"FED7", X"FE49", X"000E", X"00ED", X"FCEE", X"F790", X"FBFA", X"FBFD", X"01D4", X"FEAC", X"FFB0", X"034F", X"02D2", X"061B", X"0209", X"025A", X"016D", X"0208", X"00DC", X"01D3", X"FF1F", X"FD75", X"0335", X"0405", X"039C", X"044C", X"01E1", X"0221", X"0222", X"015B", X"0182", X"FF14", X"FA37", X"FA7D", X"FC9D", X"FB5B", X"FCDF", X"FE6D", X"037D", X"01DB", X"0412", X"0692", X"0469", X"0474", X"0246", X"01B6", X"0020", X"FFB9", X"FF8C", X"FF68", X"0354", X"0328", X"03F0", X"048A", X"02FF", X"0284", X"0400", X"0608", X"04EE", X"01F3", X"FD51", X"F962", X"FB61", X"FBE5", X"FE26", X"FEFB", X"018D", X"010B", X"00B7", X"046C", X"0665", X"03C0", X"02E0", X"02A1", X"009D", X"0113", X"01D5", X"0133", X"0147", X"0058", X"0431", X"0449", X"038B", X"03F9", X"0441", X"0680", X"04AF", X"0566", X"FD22", X"F705", X"F900", X"0175", X"FF67", X"010A", X"027E", X"035A", X"FFAE", X"00C1", X"0255", X"026C", X"01B0", X"FFC2", X"FF8F", X"FF8A", X"0215", X"01CB", X"FE72", X"FF2C", X"0200", X"0142", X"02B8", X"032F", X"02BE", X"0200", X"04AF", X"00E1", X"FCF3", X"FA53", X"F6C0", X"FCAA", X"FE09", X"003C", X"02EB", X"024F", X"FF61", X"002D", X"FF1F", X"FDDB", X"FDD2", X"FD32", X"FD1A", X"FD71", X"FEA4", X"FDE1", X"FC3D", X"FE29", X"005E", X"FF61", X"0234", X"001E", X"0034", X"01CC", X"0257", X"0047", X"FD58", X"FAF4", X"FBA9", X"FEF8", X"FC22", X"038D", X"00C1", X"030D", X"0369", X"0090", X"FD08", X"FBD5", X"FA10", X"F826", X"F87D", X"F9D6", X"FC11", X"F973", X"FA4B", X"FBC2", X"FDAD", X"FF4C", X"FF59", X"FFA8", X"FF8C", X"0060", X"017E", X"FDE9", X"FBEA", X"F7C8", X"FBD8", X"0112", X"FFA5", X"FF3E", X"FFAF", X"03D5", X"0452", X"00E4", X"FBFF", X"F864", X"F701", X"F600", X"F7DE", X"F768", X"F834", X"F75C", X"F84D", X"FB11", X"FAA3", X"FC21", X"FCFF", X"FC7F", X"003C", X"FF53", X"FDCF", X"FD13", X"FA71", X"F9FE", X"FC0C", X"FFB4", X"FE80", X"004D", X"FDA8", X"044D", X"054A", X"008F", X"FB29", X"F83C", X"F73F", X"F8CF", X"F841", X"F7B8", X"F6F0", X"F73F", X"F81D", X"FA19", X"FB43", X"FB6A", X"FBE3", X"FBA6", X"FE1A", X"FE2B", X"FC95", X"FE89", X"FC59", X"FDEE", X"011F", X"FE58", X"FE9A", X"FF63", X"0100", X"03D8", X"0571", X"0064", X"FA94", X"F955", X"FA6B", X"FA78", X"FC3F", X"FCFF", X"FA0E", X"FBC9", X"F953", X"FA56", X"FBEC", X"FD66", X"FAE2", X"FB81", X"FD72", X"FEE0", X"FC2D", X"FB62", X"FEF9", X"FE23", X"FE2A", X"FBB5", X"003B", X"FF47", X"0139", X"03DA", X"04C1", X"02BB", X"000D", X"FF77", X"0027", X"FF6D", X"FEB0", X"FFBC", X"FED1", X"FE4C", X"FEEE", X"FB31", X"FC79", X"FC31", X"FA77", X"FBF3", X"FBCD", X"FBC2", X"FD69", X"FE5D", X"FDF0", X"FEB8", X"FDEE", X"FDB8", X"FFBD", X"FFD8", X"001D", X"0297", X"072B", X"0657", X"049B", X"0748", X"041D", X"0168", X"004E", X"007D", X"FFC9", X"FD65", X"FDE6", X"FD6F", X"FBA7", X"FA62", X"FC80", X"FC1E", X"FC6D", X"FCD3", X"FF9C", X"FF73", X"FF34", X"0044", X"FDED", X"FFA0", X"0016", X"FF4D", X"0084", X"020A", X"05CE", X"0A0E", X"0831", X"0A24", X"09E4", X"051F", X"0284", X"0470", X"010F", X"FF0C", X"FE35", X"FE49", X"FD78", X"FD10", X"0190", X"FCB5", X"FB6D", X"0219", X"04AF", X"0485", X"02C2", X"FEB5", X"FCBB", X"FE29", X"001B", X"FF1D", X"FFDB", X"00E6", X"0402", X"0776", X"0955", X"075F", X"0705", X"0673", X"04B9", X"02CD", X"02DC", X"0311", X"0144", X"0158", X"FF7D", X"0047", X"0040", X"0061", X"03A4", X"0671", X"073D", X"0514", X"03BA", X"0164", X"005E", X"FDCE", X"00D2", X"FF1F", X"0019", X"002C", X"FF10", X"00AF", X"0439", X"057B", X"04DA", X"04EF", X"0635", X"053A", X"00DA", X"0219", X"0555", X"0843", X"09AF", X"0818", X"03B4", X"0404", X"054A", X"04EA", X"066F", X"03F7", X"FFA3", X"0014", X"0016", X"FDB1", X"FFF9", X"0062", X"0091", X"001A", X"00B1", X"0126", X"013E", X"021D", X"01CD", X"0317", X"02DB", X"049A", X"FE79", X"FF54", X"02F2", X"0496", X"0307", X"01F6", X"0447", X"02F0", X"00F8", X"02CE", X"03BA", X"0371", X"02FD", X"005B", X"01AE", X"FFCC", X"019A"),
--        (X"FF9F", X"0018", X"FF91", X"FEC0", X"FF77", X"00C1", X"FF19", X"00FD", X"FF92", X"FF8B", X"0060", X"00B8", X"0084", X"0078", X"FD98", X"0060", X"00AE", X"00C3", X"FF76", X"FF63", X"00B6", X"FFDE", X"0073", X"FFBF", X"FE43", X"0072", X"FFBD", X"00C2", X"FF89", X"0001", X"010D", X"01ED", X"FFA1", X"0011", X"FF2D", X"FFEC", X"FFEF", X"020B", X"00B4", X"011E", X"0359", X"01B0", X"01D9", X"FFB9", X"FB70", X"FCE7", X"02D2", X"032A", X"0262", X"00F2", X"00B1", X"001D", X"00E8", X"00D0", X"0060", X"FFB4", X"FF85", X"FF66", X"FF9E", X"FDE5", X"00D4", X"032C", X"020C", X"015E", X"0149", X"FF73", X"FF7B", X"FFEB", X"FFDF", X"FF31", X"037E", X"04AC", X"022E", X"02DD", X"0570", X"06B2", X"050F", X"031C", X"0368", X"FFEE", X"FDC3", X"FD93", X"00DD", X"0092", X"FF09", X"00A1", X"00A6", X"FF55", X"01AD", X"0032", X"00BB", X"FDC0", X"FD5B", X"FCD9", X"FB8C", X"F92D", X"F9BE", X"FB6B", X"FD20", X"0095", X"0097", X"028E", X"0542", X"07FD", X"03FE", X"0781", X"077E", X"0504", X"FFAD", X"FD86", X"FEF6", X"FFBD", X"009A", X"FF67", X"00E7", X"FDDB", X"0109", X"00A1", X"FD6E", X"FCFC", X"FAE6", X"F9E4", X"F86B", X"F806", X"FA88", X"FB4C", X"FD84", X"FEB4", X"0347", X"024F", X"06A0", X"06F1", X"082E", X"09A8", X"0874", X"089F", X"06C2", X"0321", X"0154", X"00D8", X"FF93", X"FFFF", X"FF13", X"FD2A", X"FF6D", X"FE43", X"FDCB", X"FD11", X"FB58", X"FC1E", X"FC1C", X"F98F", X"FB51", X"FB3B", X"FEC8", X"011B", X"00DF", X"015D", X"02E1", X"032A", X"0553", X"065A", X"091A", X"0AC9", X"0977", X"0263", X"0411", X"0214", X"0113", X"FECD", X"FD61", X"FB57", X"FF3C", X"FF76", X"FE9F", X"FFC5", X"FE1B", X"FE08", X"FBF8", X"FB27", X"FAC6", X"F831", X"F8F9", X"FACA", X"FA8D", X"F95F", X"FB95", X"FD8B", X"FFC5", X"FFB4", X"04B7", X"0AA7", X"0932", X"05D3", X"03B8", X"0043", X"FFA1", X"FE2F", X"FD03", X"FAD5", X"FEB0", X"0188", X"0025", X"0247", X"FCE0", X"FE0E", X"FAEB", X"FB12", X"F7EF", X"F8A0", X"F806", X"F738", X"F742", X"F7FA", X"F8EF", X"FA6A", X"FA06", X"FC32", X"0096", X"0613", X"07F2", X"05D2", X"0466", X"010D", X"FEE5", X"FDC3", X"FD69", X"FE52", X"FDEA", X"013F", X"FED7", X"009D", X"FD81", X"FDE0", X"FB5F", X"FC6E", X"FA1E", X"F7D0", X"F3D1", X"F3E6", X"F4D8", X"F89B", X"F954", X"F897", X"FACB", X"FC5A", X"FCBA", X"0053", X"060F", X"0611", X"01F3", X"0123", X"FFC3", X"0091", X"FFE1", X"FB4B", X"0042", X"FFBA", X"0159", X"FF36", X"0190", X"FFB6", X"FE16", X"00D9", X"FD26", X"FBC1", X"F688", X"F7F7", X"FA13", X"FAE1", X"FAFD", X"FC2E", X"FCE1", X"FD5B", X"FD28", X"FE5B", X"035C", X"065C", X"03F5", X"004D", X"FF01", X"FFE4", X"FE76", X"FCF2", X"0406", X"023F", X"0227", X"032A", X"029F", X"0278", X"02C1", X"0247", X"0342", X"01C4", X"FF5D", X"006F", X"00A4", X"FE3E", X"FF03", X"FF27", X"FDF9", X"FCD7", X"FB77", X"FDB7", X"0294", X"0561", X"02E6", X"FF08", X"00A9", X"0023", X"FF18", X"00B0", X"03D3", X"03E9", X"03DC", X"03AB", X"028F", X"0403", X"0469", X"0443", X"04D0", X"0515", X"0370", X"0486", X"03CF", X"FFEE", X"FEF2", X"FE65", X"FC9B", X"FB4E", X"FB21", X"FF7F", X"FF26", X"012E", X"FF84", X"0012", X"FFC3", X"0010", X"01BE", X"03CF", X"0097", X"0516", X"04E1", X"0622", X"0409", X"02F2", X"0433", X"0540", X"07A0", X"044B", X"0376", X"043D", X"01E1", X"003E", X"FFEA", X"FDBD", X"FE32", X"FD33", X"FF38", X"00E4", X"0167", X"0158", X"FF80", X"FF1D", X"00AB", X"000F", X"0158", X"02FD", X"0108", X"03F5", X"0653", X"0570", X"031C", X"0381", X"021E", X"034E", X"02DF", X"019B", X"0238", X"0320", X"00AD", X"015C", X"00B3", X"0175", X"00C3", X"0093", X"03F3", X"0357", X"045A", X"000C", X"FC73", X"FCED", X"019B", X"001E", X"015D", X"0367", X"00FA", X"056D", X"0377", X"0104", X"029B", X"02B3", X"FFD6", X"001A", X"FFA4", X"00D4", X"03DD", X"02B8", X"0131", X"0009", X"00C7", X"01C7", X"00AA", X"018B", X"039E", X"05AE", X"03F0", X"FE8E", X"F784", X"FF17", X"00E3", X"01CD", X"02AD", X"0417", X"FDA7", X"FF19", X"012C", X"0121", X"0285", X"0034", X"FEB5", X"FEDD", X"012B", X"0487", X"05F3", X"03BA", X"0084", X"FEBC", X"00A4", X"0296", X"00BC", X"00D3", X"02D8", X"0290", X"00C7", X"FE0D", X"F771", X"FB24", X"FF21", X"FF95", X"FF1D", X"FEB0", X"F8CF", X"FCE2", X"FFEA", X"FF80", X"0064", X"FD3F", X"FC37", X"FFCF", X"0037", X"053A", X"0714", X"0323", X"004D", X"0037", X"003A", X"01EB", X"0218", X"00A1", X"01B5", X"0240", X"FDF2", X"FA10", X"F8BA", X"FC12", X"FF7D", X"0058", X"FD5C", X"FBDA", X"F994", X"FE66", X"FF4F", X"FEEC", X"FE11", X"FE03", X"FF7A", X"0088", X"01CF", X"0592", X"0724", X"0241", X"0108", X"0017", X"FFFC", X"0105", X"01C1", X"011D", X"FCCC", X"009B", X"FDC3", X"F940", X"F9CC", X"FC6A", X"FD8C", X"FF17", X"FD17", X"FAA6", X"FAF7", X"FEA1", X"FE25", X"FD63", X"FE91", X"FF6C", X"FF8C", X"00CE", X"02AD", X"053E", X"042C", X"01E9", X"0279", X"000F", X"FF37", X"00E0", X"00BC", X"0039", X"FD0B", X"FBE7", X"FB8B", X"F988", X"FD59", X"0049", X"016F", X"007F", X"0157", X"FC91", X"F9E8", X"FDBA", X"FD64", X"FEC2", X"FF0F", X"FF0A", X"FFBC", X"0243", X"025E", X"01D8", X"030C", X"016C", X"00D8", X"0128", X"FF6B", X"FE1E", X"FE0A", X"FFC6", X"FD1A", X"FD82", X"FDDD", X"F963", X"FC95", X"013E", X"FFC9", X"FDB5", X"FF8E", X"FC8A", X"FAD9", X"F7F3", X"FCFE", X"FD71", X"0080", X"0091", X"02DA", X"02F5", X"0322", X"022B", X"01A3", X"0363", X"0149", X"022A", X"02B3", X"FEE4", X"FDA7", X"FDD6", X"FD76", X"FFBA", X"FDC9", X"FA95", X"FF14", X"FF66", X"001E", X"FF2A", X"FBC9", X"00DD", X"FEA1", X"FD52", X"FB1D", X"FD99", X"0064", X"0067", X"0066", X"01FB", X"0238", X"02DC", X"0420", X"037D", X"00DA", X"0465", X"0149", X"00D4", X"033C", X"0144", X"00FE", X"FCEE", X"FDCD", X"FD32", X"00B8", X"00FF", X"0081", X"FFBD", X"FAFE", X"FDB6", X"0065", X"FEDE", X"FBF4", X"FD06", X"FD5E", X"FEC6", X"FFC5", X"FFEB", X"FED7", X"0068", X"015F", X"02FF", X"0265", X"045B", X"02C4", X"01CD", X"FFEA", X"00B9", X"FD7F", X"FC27", X"FDD4", X"0053", X"03F4", X"FF42", X"0055", X"0058", X"FC84", X"FB19", X"0110", X"FF2A", X"FFB4", X"FC40", X"FCAB", X"002C", X"FE31", X"FE45", X"FF2E", X"FEDC", X"0185", X"015A", X"021B", X"026A", X"025C", X"FF5B", X"0176", X"FBB3", X"FC6C", X"FC69", X"FC13", X"0095", X"049A", X"FF7C", X"FF82", X"00A9", X"009F", X"FC19", X"FBB7", X"FDCE", X"FCED", X"F9BE", X"F8ED", X"FE27", X"FE1D", X"FE24", X"FE9B", X"FCA1", X"FEAE", X"FB27", X"FC74", X"FC0A", X"FE9F", X"FD72", X"FD8E", X"FD6B", X"FC3D", X"FBED", X"FC6C", X"0141", X"02D9", X"FFCB", X"FE8E", X"00E5", X"014B", X"007F", X"FB24", X"F753", X"F6D6", X"F77F", X"F57D", X"F7DD", X"F83E", X"F8ED", X"F839", X"F7F1", X"FA4E", X"F8A0", X"F7E3", X"F8CF", X"F756", X"F674", X"F824", X"F94E", X"FBE6", X"FEA9", X"FFE7", X"FE65", X"FFF8", X"FF43", X"FFCC", X"00D1", X"0066", X"FCE6", X"FB90", X"F99E", X"F74C", X"F6D9", X"F479", X"F2F0", X"F375", X"F5B1", X"F35B", X"F216", X"ED7B", X"F30E", X"F305", X"F338", X"F039", X"F4DF", X"F748", X"F99A", X"FD7B", X"FE4B", X"FDD4", X"0033", X"FFB9", X"002D", X"0153", X"FFEC", X"FFF5", X"015A", X"0078", X"0146", X"FECF", X"FE66", X"FC68", X"FB2E", X"F9BB", X"FC1D", X"FAD9", X"FD29", X"F78A", X"F89F", X"F8D9", X"FAAF", X"F936", X"FCB2", X"0177", X"FFF2", X"009E", X"0118", X"FF43", X"FEB8", X"0074", X"FFF2"),
--        (X"001B", X"FEF3", X"00F8", X"FFF5", X"FFB3", X"FFBD", X"0024", X"FFD6", X"007B", X"0112", X"FFCB", X"00EB", X"0100", X"0085", X"0045", X"00F0", X"00CF", X"FFDF", X"FF50", X"0076", X"0040", X"FFE6", X"FF25", X"0186", X"FF1D", X"FFDB", X"0062", X"0054", X"FFFD", X"0107", X"FF6D", X"FFD9", X"00C1", X"00AE", X"FF7A", X"FF13", X"FEB7", X"012E", X"FFC3", X"FE17", X"FC7F", X"FD42", X"FE0B", X"FFE3", X"021C", X"FF6F", X"FCF5", X"FBEB", X"FD7D", X"FE3F", X"002B", X"FFA4", X"008C", X"00CF", X"00E2", X"FF8A", X"0024", X"FF3A", X"FF9A", X"FE7E", X"FDEE", X"FF36", X"0029", X"FF9E", X"0001", X"009E", X"FCDA", X"FD11", X"FE04", X"FDCA", X"FCD3", X"FE87", X"FE65", X"FF18", X"FBEC", X"F9F3", X"FABC", X"FB4B", X"FB15", X"FBAC", X"0010", X"021C", X"018E", X"0053", X"00DA", X"00FD", X"00C9", X"FFBB", X"FF96", X"FCA6", X"FECF", X"FEED", X"00CA", X"03C4", X"003F", X"FF52", X"FFAF", X"FE89", X"FB00", X"FB81", X"FBC0", X"F9AF", X"FCF9", X"FAA0", X"FBC2", X"FDFB", X"00C1", X"FB94", X"FBDF", X"FFAB", X"FCC8", X"FE7F", X"00B6", X"0062", X"020F", X"FD31", X"FC66", X"FE81", X"FEEB", X"FEA6", X"00A7", X"0118", X"FFDF", X"FF2C", X"003D", X"FE75", X"00E8", X"0066", X"0095", X"0171", X"FE93", X"FDC8", X"00C6", X"FFCD", X"FE39", X"FFF5", X"0139", X"0178", X"0465", X"00D6", X"FF2C", X"001F", X"01CF", X"FB72", X"FD27", X"00AF", X"FF84", X"FFD4", X"025F", X"022A", X"011D", X"00BF", X"018B", X"0047", X"0024", X"FEA7", X"FF52", X"FF55", X"FD6C", X"FD94", X"FFFC", X"02DF", X"0273", X"0175", X"02CD", X"0418", X"03EA", X"0019", X"0007", X"FF26", X"0231", X"FFB6", X"0298", X"03D4", X"01B5", X"031C", X"01FA", X"0113", X"003A", X"0165", X"0133", X"FD2D", X"FDB3", X"FD76", X"FDDB", X"FC7E", X"FE27", X"FF99", X"0097", X"0323", X"0119", X"0108", X"03AC", X"03D2", X"0349", X"0315", X"FF6D", X"0174", X"03BA", X"FEF2", X"FFEC", X"03C4", X"0334", X"03DD", X"0348", X"02A0", X"00B2", X"00BF", X"FFBC", X"FE51", X"FD16", X"FD5C", X"FF13", X"FE21", X"0048", X"017D", X"0254", X"030D", X"0511", X"052A", X"04D0", X"02D3", X"0203", X"04DE", X"FE4C", X"037D", X"03D3", X"FFE8", X"0042", X"0236", X"0341", X"0429", X"028A", X"02FC", X"027E", X"039D", X"01C2", X"0276", X"0012", X"FFB2", X"0087", X"0097", X"0068", X"025D", X"0213", X"0207", X"02A9", X"063B", X"05DD", X"049B", X"0306", X"02CC", X"01D4", X"02C8", X"029E", X"0238", X"0386", X"04A9", X"031E", X"0381", X"0389", X"03C6", X"0313", X"0572", X"04B2", X"03A8", X"02CB", X"022B", X"00C8", X"02F8", X"012B", X"01E0", X"0016", X"018A", X"026D", X"0363", X"06C7", X"092A", X"0719", X"018B", X"021C", X"0516", X"00D4", X"FCFF", X"02CC", X"056E", X"0417", X"039A", X"046C", X"04C1", X"0544", X"04C6", X"04FE", X"060B", X"03E6", X"02C9", X"01B0", X"FEC4", X"FE75", X"FF44", X"FF72", X"0096", X"FF9C", X"01F8", X"04D3", X"06F1", X"0857", X"02B8", X"0167", X"01CB", X"0069", X"FB4B", X"0253", X"04D4", X"0102", X"05B6", X"028F", X"0299", X"00B8", X"FF8E", X"FD3D", X"FF35", X"FFFC", X"FDF2", X"FDA7", X"FB20", X"FC68", X"FD32", X"FC3E", X"FDBD", X"FEA4", X"FD9C", X"02F6", X"0539", X"0627", X"0228", X"0186", X"0241", X"025A", X"FB7F", X"00F7", X"00A5", X"FF56", X"00AC", X"0294", X"FF59", X"FC7C", X"F940", X"F69B", X"F980", X"FA60", X"FA29", X"FABE", X"FA54", X"FB36", X"FB92", X"FC2E", X"FC84", X"FB40", X"FAE2", X"FE06", X"07D9", X"06BF", X"02F5", X"00C5", X"01F7", X"0458", X"FB05", X"F99C", X"F956", X"F9C1", X"FB8D", X"FB93", X"FC20", X"F9AB", X"F6E0", X"F6F7", X"F9AC", X"FA3B", X"FBC2", X"FA52", X"FAC6", X"FA55", X"FB71", X"FCC6", X"FC4E", X"FAFD", X"F9CE", X"FC60", X"03ED", X"088E", X"042E", X"0077", X"FE20", X"FE8A", X"F98F", X"F5EC", X"F634", X"F67A", X"F658", X"F74F", X"F74B", X"F828", X"F7AE", X"F777", X"0135", X"FD53", X"FDF6", X"F941", X"FBB1", X"FD6E", X"FC7B", X"FD81", X"FDD6", X"FD33", X"F970", X"FC43", X"040E", X"084B", X"02F8", X"0202", X"FCA2", X"FE33", X"FAE7", X"F6D3", X"F39B", X"F4DC", X"F40B", X"F3F7", X"F7A5", X"F7A5", X"F9A0", X"FFC6", X"0361", X"0228", X"FFA0", X"FE49", X"FD1D", X"FD7E", X"FAC6", X"FB45", X"FECD", X"FD98", X"FCE4", X"FEE3", X"0502", X"0C49", X"0395", X"00B3", X"FAA8", X"FD0D", X"FDD0", X"F80D", X"F530", X"F518", X"F374", X"F6C0", X"FA09", X"FC2D", X"007F", X"01C7", X"0345", X"0246", X"03BE", X"01F5", X"FFD5", X"FD5B", X"FB5B", X"FDCE", X"FDBA", X"FEE5", X"FD72", X"00F5", X"072B", X"09D3", X"03D0", X"0082", X"FDEC", X"FC4D", X"FF91", X"FAE8", X"F8AB", X"F9AE", X"F9F7", X"FA6D", X"FE34", X"0168", X"0318", X"0528", X"03DF", X"037D", X"0255", X"0069", X"FDE2", X"FD8F", X"FD2D", X"FBDB", X"0007", X"FD65", X"FC78", X"00FC", X"06B9", X"073F", X"04DA", X"0269", X"FF5B", X"FD07", X"FF19", X"FE84", X"FADD", X"FC70", X"FDE9", X"FF31", X"0104", X"0290", X"052E", X"0502", X"047B", X"0336", X"0391", X"0079", X"FFEC", X"FE69", X"FD14", X"FDA2", X"FD1E", X"FD4E", X"FE9B", X"01F1", X"04E3", X"058B", X"03CC", X"FF74", X"0037", X"FF9B", X"FDFA", X"FEBF", X"FD40", X"FEBE", X"FFE5", X"023C", X"0514", X"04A9", X"01F6", X"0379", X"0572", X"03BE", X"0230", X"004D", X"0124", X"FFCA", X"FDF2", X"FF1D", X"FDB5", X"FC38", X"FE33", X"FFF2", X"06FB", X"04DF", X"036E", X"FF66", X"FEC9", X"FFDE", X"FBF8", X"FDD3", X"FF3E", X"00E6", X"00E0", X"029B", X"038F", X"047B", X"0409", X"0566", X"0258", X"00FA", X"01A6", X"028B", X"FF89", X"FF0C", X"00BA", X"FE09", X"FEE8", X"FF19", X"FEC6", X"015B", X"029B", X"0368", X"FEDD", X"FF35", X"0054", X"FCC7", X"FDBF", X"FC41", X"FFFD", X"0112", X"0206", X"01C0", X"0185", X"03A3", X"0259", X"00B4", X"020E", X"0055", X"00F7", X"0116", X"02C0", X"013F", X"006A", X"0081", X"FFE6", X"FE69", X"0042", X"0392", X"04F5", X"006B", X"FE74", X"FF7E", X"FF74", X"FD38", X"FCDA", X"FEB8", X"FE96", X"0226", X"0150", X"016E", X"013B", X"007C", X"0196", X"01AA", X"013F", X"023F", X"FFCC", X"0101", X"FFB2", X"FF4C", X"FEA5", X"0001", X"0327", X"FFC4", X"0004", X"037D", X"0299", X"FD76", X"FF21", X"FDDC", X"00EF", X"FFE9", X"FA09", X"FB8E", X"FBA0", X"FECE", X"FE5D", X"FF57", X"0183", X"FF9F", X"003E", X"03AF", X"01CE", X"0367", X"0297", X"0101", X"0001", X"0071", X"01CD", X"02E6", X"0178", X"0134", X"FFC2", X"FE12", X"0146", X"0062", X"00A9", X"0059", X"008F", X"001E", X"F8FA", X"F877", X"F978", X"F88E", X"FACD", X"FD52", X"FED3", X"FE9D", X"0096", X"007D", X"02FA", X"0253", X"021C", X"FFE8", X"01B0", X"041B", X"0412", X"0317", X"FEBF", X"FBF3", X"FBB6", X"040C", X"0254", X"0367", X"FFDC", X"0110", X"0074", X"FE5B", X"021E", X"FC26", X"FA06", X"F974", X"FA8A", X"FB09", X"FD13", X"FC4A", X"FE87", X"0122", X"FF69", X"015C", X"00BF", X"0266", X"027E", X"03EC", X"FFAB", X"FD4A", X"FC73", X"FCF4", X"FD43", X"FF25", X"00D1", X"026C", X"0092", X"0084", X"FF45", X"0047", X"0084", X"FE6F", X"FBEE", X"FDAD", X"004C", X"0325", X"020C", X"00FD", X"03AC", X"FF50", X"FDD5", X"FCC7", X"FE3C", X"FE72", X"FFBF", X"FDD7", X"FCF3", X"FA81", X"FBE9", X"FEB2", X"FFA5", X"0014", X"FF76", X"FFD8", X"FDC5", X"FF6F", X"00E8", X"FFA3", X"FFD0", X"01E8", X"01C6", X"02A0", X"0220", X"06B6", X"0441", X"079E", X"0167", X"02D9", X"0904", X"0418", X"01F5", X"066D", X"05D8", X"0140", X"03DB", X"FEFF", X"FE5A", X"FD88", X"0397", X"FFEE", X"00AE", X"0170", X"FF95"),
--        (X"FE61", X"FFC2", X"0050", X"0009", X"FF6F", X"0003", X"005F", X"FF81", X"FFA4", X"FF22", X"FF9D", X"0077", X"00F6", X"0014", X"FFA2", X"FEF4", X"FF0B", X"00A5", X"00F1", X"FF08", X"0052", X"FFEB", X"FEC1", X"0131", X"FEF2", X"00E6", X"FF51", X"017B", X"0058", X"001D", X"FFF8", X"FEF8", X"FFB7", X"FFC6", X"FEF7", X"00FB", X"00E8", X"000C", X"FFAB", X"0089", X"02AB", X"033F", X"FF77", X"FF09", X"01D8", X"0144", X"FFA0", X"FEF2", X"FEC0", X"FE4F", X"FEBC", X"0085", X"FF63", X"0053", X"FF99", X"FF6F", X"FE29", X"FFC8", X"0025", X"FE44", X"0108", X"0127", X"023C", X"01EA", X"0344", X"048B", X"03AC", X"03DD", X"039A", X"02EB", X"018F", X"0135", X"043B", X"0680", X"0641", X"056E", X"02A3", X"018A", X"002E", X"00BE", X"0204", X"0015", X"00BF", X"FF2C", X"0076", X"FF9B", X"FF17", X"FD3D", X"013D", X"00CC", X"0116", X"012C", X"FF7B", X"02FF", X"00A3", X"FE07", X"FCEC", X"FE13", X"FD9F", X"FC4E", X"FD37", X"FDB7", X"FD5C", X"006C", X"010E", X"03D2", X"0303", X"046F", X"0392", X"004E", X"02B2", X"FF1E", X"0021", X"FF22", X"FCE3", X"FC49", X"FEA0", X"0074", X"FF7E", X"FFF8", X"FE49", X"00C5", X"FE2A", X"FE6B", X"FC83", X"FBC4", X"FC16", X"FDE4", X"FF02", X"0137", X"0025", X"FF13", X"0090", X"01A0", X"021C", X"050A", X"0303", X"FE0D", X"FE0D", X"00C4", X"FFD6", X"FF3B", X"FFC4", X"FFF2", X"FFB6", X"FC8E", X"FE26", X"000D", X"01D1", X"02E5", X"00E1", X"0096", X"FFB0", X"FE57", X"FF19", X"FFD2", X"0014", X"01D9", X"0317", X"FFD2", X"036C", X"0201", X"03A1", X"05E5", X"021A", X"0095", X"FF6B", X"0183", X"0150", X"001A", X"FB42", X"FC2D", X"FF4A", X"FE48", X"FFCC", X"0250", X"00EB", X"00A0", X"FF4F", X"FE0B", X"FE96", X"FC54", X"FDCF", X"FD83", X"FD8E", X"FD83", X"FC8C", X"00F1", X"FF8D", X"015D", X"04A9", X"0599", X"04CE", X"00B6", X"018C", X"01DB", X"00CE", X"FC6A", X"FEE1", X"F99C", X"FE28", X"00D7", X"014B", X"02F1", X"0137", X"0028", X"FF71", X"00C3", X"FDE5", X"FF1D", X"FCE2", X"FC11", X"FD3C", X"FD73", X"FBDC", X"FB2B", X"FD43", X"FF85", X"032C", X"03D7", X"0830", X"03DD", X"006A", X"02D6", X"041C", X"FF51", X"FF57", X"F9E1", X"FB4A", X"0141", X"009B", X"029F", X"00FD", X"01FE", X"0002", X"024A", X"FF60", X"FE84", X"FE2C", X"FE05", X"FD78", X"FCC3", X"FAEA", X"FB45", X"FE0E", X"FD5E", X"FFF5", X"06C9", X"0A12", X"060D", X"0179", X"FF47", X"FEF7", X"FD34", X"FFB9", X"F9FC", X"FD4E", X"0071", X"FFFC", X"00B8", X"000A", X"01B7", X"0348", X"04BE", X"0281", X"0041", X"FBB5", X"FCD5", X"FDE0", X"FD3E", X"FC0F", X"FCDA", X"FB5E", X"FE3C", X"FF1E", X"06C8", X"0B49", X"0958", X"03AB", X"FCE7", X"FF3B", X"FDEE", X"FABE", X"FB4B", X"FF83", X"00D6", X"FD52", X"FD91", X"FFA2", X"0194", X"0456", X"04AF", X"0610", X"FE6C", X"FCB8", X"FD56", X"FC58", X"FCB3", X"FBE9", X"FB68", X"F9C6", X"FA73", X"FC3D", X"05A7", X"0E11", X"0A4B", X"0535", X"FDEC", X"00AD", X"FE34", X"FC04", X"FBD5", X"FFA4", X"FFD0", X"FF89", X"FD88", X"FE4E", X"011A", X"FFE5", X"0286", X"0211", X"FAF1", X"F8C4", X"FBE8", X"FF20", X"FA6A", X"F955", X"F98C", X"F8C1", X"F95F", X"FA3C", X"00A9", X"0B08", X"093B", X"03D8", X"FCAD", X"00AF", X"00A6", X"FDF1", X"FBCA", X"FE36", X"FDF6", X"FD1F", X"FC9D", X"FE03", X"FEC0", X"0253", X"049E", X"04A3", X"FA30", X"F930", X"FA54", X"FC0C", X"FB96", X"FB98", X"FBAD", X"F9B7", X"FA92", X"FBEC", X"FE7E", X"0401", X"02F2", X"029F", X"FD8A", X"FFD4", X"00CF", X"FFC8", X"FC73", X"FB97", X"FFFF", X"FFA6", X"FFB5", X"FFD1", X"0067", X"02D6", X"05FD", X"0515", X"FC54", X"FA94", X"FC27", X"FAE6", X"FDF0", X"FE36", X"FFFF", X"000D", X"FF48", X"0487", X"05B3", X"05E1", X"02E5", X"03AF", X"0378", X"01F7", X"0001", X"FDBB", X"FD26", X"FFD3", X"010A", X"00BD", X"019E", X"0155", X"0229", X"0515", X"0735", X"0555", X"FCDC", X"FB67", X"FDE6", X"FFDC", X"0206", X"0006", X"0142", X"02A5", X"00E9", X"0354", X"0391", X"0711", X"0623", X"04E6", X"00C2", X"0241", X"FD4D", X"01CD", X"FFC5", X"0027", X"0151", X"0074", X"014C", X"014E", X"0230", X"0350", X"050C", X"049E", X"FF9D", X"FDAC", X"FF99", X"015F", X"011A", X"011B", X"FFC7", X"000A", X"018E", X"006B", X"01EF", X"06AF", X"06FE", X"05AF", X"01F0", X"FDB1", X"FD02", X"FDE1", X"FEAD", X"FCC5", X"0198", X"02F5", X"0106", X"FFDE", X"00B2", X"004F", X"0382", X"0399", X"FFC7", X"FFF2", X"03BB", X"03CF", X"003A", X"FFF0", X"0056", X"0241", X"011A", X"018A", X"04F5", X"0650", X"09F9", X"041F", X"012C", X"FF83", X"FCC4", X"FFE9", X"FED5", X"FE1F", X"025F", X"056E", X"0184", X"FF46", X"FF92", X"0260", X"028C", X"014B", X"00AA", X"00C0", X"024C", X"02F0", X"FE92", X"00B9", X"FD99", X"00C7", X"027B", X"0350", X"06DD", X"096C", X"0841", X"0151", X"FF09", X"FC9B", X"0013", X"FE4E", X"FC5C", X"0056", X"039E", X"0414", X"0315", X"007C", X"003A", X"0225", X"0389", X"04EA", X"0326", X"00A8", X"0290", X"0169", X"0019", X"FE54", X"FFDD", X"004B", X"00E8", X"04B5", X"0C04", X"0BF5", X"063E", X"FF45", X"FF97", X"0091", X"FD39", X"00EC", X"FE89", X"00B2", X"029D", X"0291", X"01CD", X"027E", X"0000", X"008E", X"03DC", X"048D", X"02EC", X"0242", X"0273", X"00E2", X"FFBF", X"0108", X"003E", X"002A", X"0337", X"0734", X"0A37", X"0952", X"024A", X"00FF", X"FE69", X"0020", X"0211", X"00EF", X"FFCB", X"020C", X"01F9", X"00CA", X"FFF0", X"012D", X"00DD", X"00C9", X"04D2", X"039E", X"032D", X"0194", X"0473", X"0378", X"0231", X"025F", X"01D8", X"030E", X"0498", X"090C", X"0A64", X"0807", X"027A", X"00C4", X"000C", X"FF88", X"01A5", X"FE19", X"0209", X"03AA", X"022F", X"01B2", X"00CC", X"0150", X"0311", X"0282", X"02D4", X"044A", X"0220", X"03C8", X"024D", X"0372", X"05A9", X"01A7", X"033B", X"03B7", X"0652", X"095D", X"0D8C", X"0874", X"02E3", X"045B", X"FF8C", X"005E", X"FFF1", X"FE96", X"0224", X"022C", X"0041", X"FE5D", X"011C", X"02DC", X"02E7", X"0119", X"0012", X"01A9", X"005B", X"FDDA", X"FFAA", X"0031", X"0129", X"0253", X"023F", X"053B", X"0854", X"09CB", X"0A44", X"0869", X"0391", X"00BC", X"FFD1", X"003E", X"0021", X"FF87", X"FFA5", X"01F1", X"00AA", X"FFFA", X"0028", X"01D2", X"015E", X"019B", X"0100", X"FF59", X"FCEF", X"FD64", X"FC57", X"FE4A", X"FC8F", X"FFB2", X"022A", X"040E", X"06C5", X"05BD", X"0648", X"00A1", X"01F1", X"FD67", X"002F", X"FFC6", X"FFC6", X"FE63", X"FCBE", X"FBB2", X"FC35", X"FBA1", X"FCD1", X"FD65", X"FFC3", X"FD93", X"FF41", X"FDD7", X"FEF0", X"FDBF", X"FD8A", X"FC39", X"FBCF", X"FDF6", X"FDEA", X"FF2B", X"00AA", X"0175", X"019B", X"0478", X"02A6", X"0045", X"00D5", X"0026", X"00FF", X"FFB4", X"0107", X"FCDE", X"F7DC", X"F52F", X"F461", X"F540", X"F782", X"F855", X"F914", X"F81D", X"F9A8", X"FC48", X"FCBB", X"FC2F", X"F96B", X"F8B2", X"F5D8", X"F653", X"F7EF", X"FC1C", X"00EA", X"FFCB", X"0012", X"016A", X"FF37", X"00A7", X"004A", X"FFC4", X"FEFD", X"FE65", X"FB90", X"F891", X"F668", X"F75A", X"F567", X"F7EC", X"FAAA", X"FB1D", X"F9EA", X"F578", X"F8EB", X"F756", X"FAA2", X"F7EF", X"F8F1", X"F88C", X"F7F8", X"FA4A", X"FCE0", X"FFCF", X"FFB7", X"FFAE", X"0105", X"FF7B", X"FF95", X"FF4B", X"000F", X"009D", X"FF18", X"FDE5", X"FC56", X"FD2D", X"FC35", X"FEAA", X"001D", X"FDCB", X"FDD3", X"FA78", X"FBCC", X"FC76", X"FACC", X"F9B5", X"FB27", X"FD9E", X"FBEA", X"FC72", X"FC53", X"FF8D", X"FFC1", X"0098", X"FFB9"),
--        (X"FFB2", X"FF9F", X"00A0", X"0032", X"0158", X"011B", X"FF62", X"00CF", X"FF79", X"FF51", X"FFFD", X"FF2B", X"FEB2", X"00D3", X"001F", X"FF70", X"0023", X"001A", X"FFB7", X"00CA", X"0111", X"0035", X"FEDF", X"FFA9", X"0129", X"003E", X"003D", X"FF51", X"0174", X"0141", X"00B5", X"0096", X"0070", X"FFFB", X"01DA", X"01BC", X"018F", X"0280", X"020D", X"FDDA", X"FFDF", X"FE19", X"0058", X"FE39", X"FDB8", X"FED0", X"0078", X"01EF", X"00C4", X"00D5", X"000E", X"00F5", X"FFD3", X"00D8", X"FF70", X"00A5", X"0101", X"FDD8", X"0043", X"FF4D", X"FE4D", X"02B9", X"01FF", X"0189", X"03FB", X"02D9", X"052E", X"022E", X"00D6", X"0067", X"0329", X"0445", X"0123", X"020C", X"0392", X"0383", X"04C0", X"02BC", X"0255", X"000D", X"FFE1", X"FF30", X"01DC", X"0148", X"00A0", X"0076", X"FD91", X"FFAA", X"FFA6", X"FF86", X"023A", X"01D4", X"032B", X"04A4", X"0328", X"00DF", X"FE3F", X"00A9", X"FEFB", X"FFA8", X"FF10", X"FF81", X"0367", X"0642", X"03F1", X"04ED", X"0608", X"0822", X"037C", X"0050", X"FFE6", X"0063", X"FFFF", X"FFA8", X"FCC1", X"FE2A", X"FF2C", X"FCC8", X"FF43", X"011A", X"007C", X"0183", X"017D", X"FE89", X"00E5", X"FF8D", X"FEAF", X"FC6C", X"FF73", X"018B", X"01DC", X"01BF", X"0565", X"0366", X"0551", X"051A", X"081A", X"06A1", X"03E0", X"0325", X"FF0B", X"FF71", X"FE53", X"FC89", X"FC95", X"FB45", X"FB9E", X"FAF3", X"FDFC", X"FE89", X"FEB3", X"0090", X"0112", X"FEDB", X"FEB9", X"FAF7", X"FCC9", X"02FE", X"FF61", X"024C", X"0342", X"0324", X"01A9", X"03D6", X"0759", X"0AF9", X"05CA", X"037D", X"002E", X"001D", X"FDB6", X"FADD", X"F8BB", X"F7B9", X"F803", X"F967", X"FB45", X"FCBC", X"FCB3", X"FDE8", X"FD1C", X"FE19", X"FE06", X"FEEC", X"FF60", X"FED1", X"FF7C", X"0130", X"0100", X"FD68", X"FEFB", X"01C1", X"0646", X"0FE1", X"08A5", X"03AE", X"FFAA", X"FB83", X"FE5F", X"FA51", X"F7E3", X"F786", X"F8A8", X"FC47", X"FD22", X"FD3B", X"FC5C", X"FE4D", X"FC01", X"FDAF", X"FDFE", X"FF38", X"FE27", X"FF91", X"FD31", X"FD9B", X"FDD9", X"FE78", X"FD29", X"004A", X"0254", X"0708", X"0877", X"0213", X"FD9A", X"FCFF", X"FD9E", X"F966", X"F7C4", X"FA3F", X"FC8A", X"FE2A", X"FF50", X"FEE7", X"FE2E", X"FD72", X"FB89", X"FDFC", X"FB88", X"FC9E", X"FD30", X"FC57", X"FD14", X"FC54", X"FD5C", X"FF3B", X"FDB5", X"FD2C", X"0219", X"0676", X"097F", X"02EE", X"FFC0", X"FD23", X"FCF8", X"F75D", X"F855", X"FA7F", X"FE46", X"FE14", X"FFCA", X"FFB7", X"FF96", X"FFB8", X"FDF0", X"FBF2", X"F87D", X"F941", X"FA61", X"FB1C", X"FB79", X"FCD8", X"FD2C", X"FD4C", X"FCB2", X"0126", X"FFD2", X"0362", X"060F", X"008A", X"016B", X"FD1F", X"FAAE", X"F9D9", X"F9E8", X"FEDC", X"FF5E", X"0175", X"0132", X"023D", X"00AE", X"00FB", X"FE8D", X"F870", X"F48A", X"F446", X"F3E0", X"F700", X"FADA", X"FC8A", X"FC27", X"FF26", X"FFFC", X"028E", X"0130", X"0121", X"033E", X"015D", X"FFDB", X"FB4E", X"F880", X"FA7D", X"FED4", X"0435", X"03F4", X"02F3", X"03C0", X"034E", X"0245", X"01FD", X"FE4C", X"FA8C", X"F60A", X"F4A4", X"F6BD", X"F967", X"FC97", X"FE4D", X"FFBD", X"FFBA", X"0297", X"020D", X"0476", X"0100", X"00DA", X"0002", X"FF53", X"FB86", X"FA92", X"FD27", X"011B", X"037A", X"04B6", X"0313", X"0372", X"0380", X"0401", X"03D5", X"04B2", X"0477", X"0225", X"FF99", X"009C", X"00EC", X"003C", X"0295", X"0252", X"02E4", X"0235", X"011B", X"FEB7", X"FD16", X"FFC4", X"FE48", X"0052", X"FCEB", X"FB13", X"0013", X"0493", X"04C0", X"0574", X"056A", X"042D", X"0574", X"046A", X"079F", X"081A", X"0AF8", X"082C", X"07FD", X"049D", X"0420", X"03A8", X"01A0", X"03E4", X"0351", X"01A3", X"FF63", X"FBD9", X"FDE6", X"FE14", X"FCA5", X"0081", X"FE9A", X"FBC6", X"01EF", X"0315", X"0480", X"04BF", X"02C5", X"0365", X"0425", X"03F9", X"0679", X"05BD", X"0850", X"067F", X"0452", X"060D", X"0359", X"0020", X"FE5B", X"FEE6", X"FE45", X"FD5F", X"FB21", X"FC24", X"FC12", X"F8BE", X"0083", X"0140", X"FF48", X"FCC2", X"0064", X"FF3D", X"0138", X"0577", X"048E", X"02E7", X"013E", X"02AE", X"0203", X"0286", X"0515", X"057A", X"04FE", X"03F0", X"012E", X"FF73", X"FEAC", X"FE11", X"FB78", X"FAE1", X"F8D0", X"F9B9", X"FBC9", X"FA06", X"FDCA", X"FF8C", X"FDB5", X"FBBB", X"FF5B", X"FE98", X"03A0", X"049A", X"0135", X"0197", X"0045", X"0147", X"0253", X"03C3", X"0389", X"0485", X"04F2", X"029E", X"FFD0", X"FF3B", X"FD5B", X"FBA3", X"FBC0", X"FB88", X"F9F0", X"F9B3", X"FC92", X"F9AF", X"FC1B", X"FFCB", X"FF38", X"FE02", X"FF95", X"FCE7", X"0161", X"0496", X"0381", X"0249", X"0171", X"001B", X"03CD", X"042E", X"02E0", X"054B", X"03F8", X"01C7", X"FF1F", X"FF20", X"FF6E", X"FECB", X"FC28", X"FA0F", X"FBAA", X"FD24", X"F9AA", X"F6EF", X"FBB8", X"FF27", X"FD7D", X"FD44", X"FE8B", X"FD56", X"01BF", X"04DF", X"049C", X"00EA", X"0278", X"0238", X"036A", X"02D7", X"0307", X"02BF", X"0229", X"01C3", X"FF1E", X"FE2D", X"FEF3", X"FDE9", X"FD6C", X"FC58", X"FFE1", X"0126", X"FB4D", X"FACE", X"FC24", X"002B", X"FC3A", X"FC72", X"FC2B", X"FD3F", X"FF9B", X"0106", X"01FF", X"FFE2", X"00F4", X"0099", X"01A2", X"FFC8", X"FFF0", X"FFCE", X"0243", X"01D6", X"00C7", X"018A", X"007B", X"009E", X"FE89", X"FF12", X"0242", X"039F", X"FAF2", X"FC95", X"FC5C", X"FFA6", X"FD5B", X"FEEC", X"F8E0", X"FAF2", X"FCA4", X"FD2F", X"FEC6", X"FCD2", X"FE46", X"FDC3", X"FDB5", X"FEA3", X"FE54", X"FD80", X"0035", X"01AD", X"026A", X"0065", X"0193", X"013B", X"00C1", X"0122", X"03B2", X"054A", X"FDFF", X"FD95", X"FF60", X"FF10", X"FEAC", X"FC15", X"FA6E", X"FB0D", X"FA39", X"FB10", X"FDA7", X"FC76", X"FEEA", X"FD7C", X"FD87", X"FDF0", X"FFD0", X"FDEB", X"FF77", X"FFCB", X"0225", X"0177", X"0197", X"022F", X"0208", X"039D", X"059B", X"0430", X"FCBE", X"FC7E", X"0043", X"FF57", X"0033", X"FD43", X"FE01", X"FC30", X"F93C", X"F79F", X"FAEA", X"FDAC", X"FE47", X"FD9D", X"FE58", X"FF47", X"FDC7", X"FD56", X"FE18", X"FFC7", X"005B", X"0083", X"0298", X"03AC", X"0360", X"0440", X"076E", X"054E", X"FE55", X"FD6F", X"FF86", X"00AF", X"00AE", X"FFF2", X"FD54", X"F9C9", X"FA65", X"F7C1", X"F85C", X"FBD2", X"FDB1", X"FD94", X"FCAD", X"FEA8", X"FE73", X"FFA3", X"FD6E", X"FFE5", X"FF4C", X"024D", X"03F1", X"0752", X"07A4", X"0639", X"094D", X"02C1", X"FF37", X"FC55", X"0078", X"01C1", X"FF6D", X"FEE6", X"FE49", X"FB15", X"FA3B", X"F936", X"FC12", X"FE56", X"FDB5", X"FE89", X"FE66", X"FF76", X"FD40", X"FE52", X"FFFE", X"0037", X"FF39", X"020E", X"0555", X"09AA", X"0669", X"0481", X"0854", X"01D1", X"0122", X"FC97", X"012A", X"0122", X"00B3", X"0012", X"00D0", X"FF7C", X"FDBD", X"FF72", X"FF66", X"FC83", X"FE0E", X"FF11", X"FDE2", X"FEB8", X"FEF6", X"00C3", X"FF02", X"0071", X"FE9A", X"FEEB", X"01C0", X"05C7", X"04EE", X"017D", X"0613", X"FCC1", X"00ED", X"FE51", X"FEC9", X"FEC2", X"FFAC", X"0021", X"00D4", X"024D", X"FFE4", X"021C", X"042F", X"0366", X"00F1", X"0141", X"0242", X"03B9", X"027C", X"0176", X"006D", X"FDC0", X"FCFE", X"FA78", X"F955", X"017E", X"00DA", X"004E", X"FFE7", X"FFEF", X"0106", X"FFF6", X"00A8", X"0083", X"00E6", X"FFA3", X"00B1", X"0087", X"0034", X"0209", X"FFFB", X"FE2F", X"FF2A", X"FCB5", X"FF74", X"FF31", X"FCC5", X"FDA2", X"FF74", X"0011", X"FBAD", X"FC63", X"FC5E", X"FDBC", X"FED9", X"FDB0", X"FD00", X"FFA4", X"FFB9", X"FFA5", X"FEFA"),
--        (X"002D", X"FF77", X"0148", X"FF8F", X"FFEB", X"FF6B", X"0079", X"FF66", X"FFEB", X"0067", X"0057", X"FFE6", X"FF73", X"FEEB", X"FDF8", X"0095", X"FF9F", X"00B7", X"0060", X"0164", X"0130", X"FFBA", X"0038", X"00BB", X"0132", X"0030", X"FF51", X"002F", X"0080", X"FF3E", X"0095", X"00D3", X"0173", X"FECC", X"FE90", X"FF1E", X"FF01", X"FF04", X"FD80", X"FCA9", X"FF63", X"FF92", X"0084", X"01DD", X"FCBD", X"FD08", X"FE3C", X"0198", X"010A", X"0044", X"FE78", X"FFA0", X"FFF7", X"FEA5", X"0032", X"004F", X"FFA2", X"FF60", X"FF6F", X"00E5", X"001F", X"01C9", X"000B", X"00C0", X"FF25", X"FE15", X"FCDC", X"FAFB", X"FB50", X"FD93", X"FF4F", X"FEC4", X"FB22", X"FA00", X"FBDB", X"FE8E", X"FFAB", X"021F", X"00F7", X"FFAF", X"FEF4", X"FF75", X"FE34", X"FF58", X"FF7F", X"0008", X"00C8", X"FEEC", X"FE68", X"00B3", X"FE49", X"FDB3", X"F998", X"FA6C", X"F8B9", X"F8C7", X"F848", X"F856", X"F9DC", X"FA7C", X"F94E", X"FA9A", X"F85B", X"FABB", X"F91F", X"FDDB", X"00D4", X"0125", X"013E", X"FFB8", X"FCB4", X"0021", X"FFA6", X"0076", X"0127", X"FF85", X"FFED", X"FE96", X"FB1A", X"FCDD", X"FA8C", X"FBF8", X"FB95", X"F8FD", X"FA41", X"FC0A", X"FE6E", X"FCE6", X"FD1B", X"FECB", X"FD6D", X"FE66", X"0082", X"FF60", X"FF33", X"FE0E", X"FD57", X"FCFB", X"FED2", X"0106", X"FE3C", X"0019", X"FF9C", X"FAC8", X"FD9A", X"FB9A", X"FCC3", X"FC2F", X"FC1B", X"FCA1", X"FBD9", X"FDD9", X"FEE8", X"FCF9", X"FEDA", X"FF9B", X"FF56", X"FDB0", X"FBCB", X"FE96", X"FF12", X"FE69", X"FDEA", X"FD85", X"FA96", X"FC6B", X"FC67", X"FDEB", X"FE20", X"0038", X"FE17", X"FBC5", X"FCF9", X"FCC6", X"FBED", X"00B7", X"FD5B", X"FD77", X"FD6E", X"FE6D", X"FD4E", X"FDE5", X"FD34", X"FE4B", X"FD53", X"FD04", X"FD2F", X"FC9E", X"FE54", X"FE0A", X"FD8C", X"00A6", X"FD40", X"FC3D", X"FC02", X"FD1B", X"000B", X"FEFE", X"FFD0", X"FF02", X"FDA1", X"FE83", X"009A", X"FFCC", X"FF6F", X"FCFA", X"FDD8", X"FB7B", X"FACB", X"FAE0", X"FB1D", X"FB5A", X"FCB0", X"FB96", X"FD5A", X"FD27", X"FDC4", X"FE7C", X"FC87", X"FF84", X"FD77", X"FB29", X"FA7E", X"FC8F", X"FF55", X"0088", X"FE4B", X"FFF4", X"FE92", X"0056", X"0095", X"000C", X"FF1C", X"FF34", X"FF79", X"FD88", X"FCEA", X"FC9F", X"F98E", X"FAB5", X"FBD5", X"FD4E", X"FD48", X"FE53", X"FEF3", X"FF33", X"0035", X"FE02", X"FB33", X"F9AD", X"FB3E", X"FCED", X"013F", X"FF6F", X"FD8F", X"FF95", X"FF5F", X"001B", X"0064", X"00A6", X"FED8", X"FF3E", X"00FF", X"FFE3", X"00F4", X"FFFB", X"FF96", X"FF6B", X"00C1", X"FF85", X"FDFC", X"01D9", X"018B", X"0202", X"020F", X"FF74", X"FE09", X"FB68", X"FDB5", X"FCED", X"017B", X"0193", X"FD7A", X"FCF3", X"00DE", X"FE8A", X"012A", X"03ED", X"FF6C", X"0194", X"03F6", X"0350", X"05A5", X"0441", X"06B6", X"0804", X"03F9", X"02C4", X"03C2", X"03EB", X"040A", X"0411", X"068C", X"0522", X"0035", X"FD56", X"FB11", X"FCD6", X"0089", X"0293", X"FE81", X"0094", X"0207", X"024B", X"033D", X"0571", X"04A7", X"041A", X"0508", X"055F", X"058A", X"0765", X"0A36", X"0831", X"0766", X"031D", X"0056", X"0389", X"080B", X"09A4", X"090B", X"060D", X"05CC", X"01D2", X"FD78", X"FE0D", X"0085", X"00EB", X"0073", X"025D", X"016A", X"03F3", X"03C8", X"0412", X"0412", X"0517", X"04B8", X"040F", X"048B", X"04E8", X"0645", X"062B", X"0454", X"026E", X"FF82", X"024F", X"02B9", X"07D7", X"09B7", X"08E8", X"0861", X"04FC", X"0091", X"0049", X"00A3", X"005B", X"0213", X"03EE", X"027B", X"04EF", X"0527", X"0414", X"0379", X"02CB", X"019F", X"04DE", X"03C2", X"0392", X"0289", X"0522", X"0624", X"02CD", X"FFC6", X"00D8", X"0214", X"03CD", X"055C", X"078F", X"03BC", X"03C8", X"FC0F", X"0000", X"FED0", X"0060", X"0152", X"02F3", X"01B7", X"02F5", X"02D0", X"02A4", X"0277", X"0203", X"0347", X"048E", X"0412", X"036A", X"0302", X"037F", X"03DB", X"045B", X"02F5", X"0215", X"00BB", X"0346", X"0403", X"01E8", X"0187", X"0067", X"FA9E", X"FF5F", X"FE90", X"FF0F", X"0041", X"0115", X"00CE", X"011A", X"01A8", X"01DB", X"012B", X"01EC", X"026A", X"01D7", X"0097", X"029D", X"028D", X"0421", X"0500", X"04A8", X"01CD", X"FFE9", X"0094", X"0017", X"027E", X"0094", X"FAF1", X"FF5E", X"FAF7", X"FBB6", X"00E0", X"FE8A", X"FE27", X"FB0A", X"FDDE", X"FFD9", X"0405", X"0653", X"078D", X"0385", X"0219", X"0212", X"FF7A", X"00B4", X"0458", X"074B", X"0653", X"058C", X"01B4", X"FFAD", X"0074", X"FE4D", X"FF28", X"FD3F", X"FB8B", X"FC36", X"FAB7", X"FC0E", X"FFD6", X"FF6A", X"FD4D", X"F964", X"FBF7", X"FEC0", X"0437", X"079A", X"0A3F", X"096C", X"0593", X"02DC", X"048B", X"052B", X"067D", X"0641", X"05A9", X"019E", X"FF20", X"FF67", X"FF68", X"FFB0", X"FEB4", X"FF81", X"FE22", X"FD08", X"FD91", X"FD0D", X"000A", X"FF38", X"FF26", X"FA31", X"F938", X"FC2C", X"0139", X"0610", X"0798", X"0810", X"097D", X"091B", X"08E5", X"0718", X"07A2", X"0347", X"0055", X"FD29", X"FE99", X"FE5B", X"FE9F", X"FE0A", X"FD81", X"FE76", X"FC63", X"FC1E", X"FD3C", X"FCBE", X"FF59", X"FEB1", X"FE03", X"F886", X"FA3D", X"FD06", X"FE26", X"020D", X"0298", X"048D", X"0519", X"05E7", X"03E5", X"0352", X"FF76", X"FDE9", X"FBEA", X"FD06", X"FDF9", X"FE7D", X"FE62", X"FCC8", X"FF72", X"FEDF", X"FD05", X"FB7B", X"FA80", X"FFFA", X"FEC8", X"FEB1", X"FBDF", X"F82E", X"F97A", X"FB77", X"FCBD", X"FEDF", X"FE2E", X"FEE9", X"FEF2", X"FC40", X"FCEA", X"FDA5", X"FB19", X"FA7F", X"FA43", X"FCB3", X"FD45", X"FD30", X"FC3A", X"FD18", X"FC6B", X"FD14", X"FC5F", X"F93A", X"FD97", X"0084", X"017A", X"FE67", X"FA72", X"F6CC", X"F987", X"FC93", X"FD0D", X"FE80", X"FAFE", X"FCD9", X"FB07", X"FACC", X"F931", X"F932", X"FAD4", X"FB71", X"FBBD", X"FD1C", X"FB08", X"FC5D", X"FCCA", X"FCF0", X"FD21", X"FA4A", X"FD1E", X"FC34", X"FC16", X"FF31", X"00B9", X"FFCE", X"FAC9", X"F9FE", X"FA21", X"FCD9", X"FD82", X"FF3D", X"FCF5", X"FCB7", X"FDB1", X"FB21", X"FBF4", X"FC72", X"FDE6", X"FC8D", X"FD98", X"FD21", X"FC13", X"FC05", X"FBB7", X"FDED", X"FBAE", X"FA59", X"FCA4", X"FE41", X"FD04", X"FDBD", X"FFD0", X"0013", X"FD03", X"F906", X"F9FC", X"FAEB", X"FCFC", X"FD96", X"FCE3", X"FE03", X"FB61", X"FC54", X"FE3E", X"FCDD", X"FD40", X"FE64", X"0011", X"FECE", X"FECE", X"FF87", X"FE8F", X"FFBE", X"FB69", X"FC0A", X"FB9B", X"FADC", X"FC64", X"FFEE", X"00C5", X"FFDD", X"FF17", X"F8E4", X"FAA5", X"FBB4", X"FA80", X"FA9F", X"FB5F", X"FD07", X"FD1A", X"FDA6", X"FC68", X"FC22", X"FC5F", X"FC80", X"FD35", X"FBA4", X"FDA3", X"00C6", X"0028", X"FE6E", X"FDE9", X"FE71", X"FAD9", X"FC65", X"FF97", X"00AD", X"0095", X"FFC4", X"FE9F", X"0247", X"0016", X"FE9E", X"FC49", X"FB11", X"FA38", X"FACC", X"FAB7", X"FB9D", X"FB77", X"F9F7", X"FD32", X"FEB0", X"FAD0", X"FCC4", X"FBD8", X"FCE2", X"FFCC", X"FDBE", X"FB32", X"FD19", X"FD37", X"FF3B", X"FE59", X"FF26", X"FF9B", X"FF4A", X"FEFC", X"FF16", X"000B", X"02A4", X"0336", X"0495", X"0436", X"03D1", X"0267", X"0176", X"FE5D", X"0088", X"0294", X"FE71", X"FDBE", X"FF4E", X"FDD3", X"FD0C", X"FCDF", X"FDF4", X"FE0D", X"01BB", X"000F", X"0003", X"FF4D", X"0066", X"002E", X"FF7F", X"FFBA", X"FF0E", X"0084", X"004E", X"00B0", X"00CC", X"0179", X"01FB", X"0075", X"0032", X"FF8A", X"00BA", X"0451", X"048E", X"03FA", X"0224", X"0438", X"02D0", X"0139", X"01A3", X"0183", X"FEC3", X"0072", X"0038", X"0033", X"FEDD"),
--        (X"008E", X"004C", X"FE52", X"0138", X"FF51", X"FFBF", X"FF8D", X"FF3E", X"0074", X"FE11", X"0060", X"FED1", X"FEEB", X"FF3B", X"0085", X"00A1", X"0041", X"0089", X"00CC", X"FF49", X"011B", X"002B", X"FF8B", X"FFFA", X"FF3D", X"00AE", X"00A9", X"FF57", X"0012", X"FFDB", X"FFFB", X"00AE", X"FF07", X"0020", X"FE4C", X"FDED", X"FEBB", X"FD4B", X"FBFF", X"FC54", X"FC01", X"FCAA", X"FC55", X"FD11", X"FA34", X"FB38", X"FD3A", X"FD03", X"FB19", X"FD3E", X"FEDA", X"FD97", X"FE88", X"0045", X"0080", X"FEBC", X"FF73", X"0052", X"0079", X"FE9C", X"FE14", X"FF38", X"FE3C", X"FCF0", X"FBD7", X"FA4F", X"F95F", X"F831", X"F7E4", X"F6C0", X"F54A", X"F7A1", X"F665", X"F7CA", X"F849", X"F815", X"F9EA", X"F989", X"F991", X"FC76", X"FDCF", X"FFD2", X"00C8", X"0057", X"FEE3", X"00C5", X"025A", X"FE86", X"FF2B", X"FE51", X"FE2D", X"FDFC", X"FAC5", X"F975", X"F754", X"F8C4", X"F5E8", X"F3F6", X"F3CF", X"F322", X"F2F1", X"F6CE", X"F4D7", X"F5BA", X"FA13", X"FB85", X"FB4F", X"FAE5", X"FAB8", X"FBF6", X"FDF8", X"0036", X"FF7F", X"FE35", X"0267", X"012A", X"00C2", X"FDBA", X"00F6", X"FF74", X"FC63", X"FCFB", X"FEDB", X"FD64", X"FB59", X"FCD7", X"FAE8", X"FBC3", X"FB8E", X"FB20", X"FB2A", X"FF32", X"FFDA", X"00F0", X"0171", X"008C", X"FA22", X"F9E3", X"FA68", X"FC61", X"0148", X"0029", X"0165", X"001D", X"0148", X"0096", X"0049", X"FE78", X"FF59", X"FE93", X"FEF2", X"01B5", X"012F", X"0030", X"000C", X"FE6C", X"FB90", X"FA25", X"F944", X"FAF5", X"FC23", X"FE3D", X"00BF", X"028F", X"FFAB", X"F906", X"FB66", X"FDF7", X"009E", X"FEF1", X"FD13", X"FD49", X"00CC", X"FEEE", X"FDE8", X"FCCE", X"FB9E", X"FFE9", X"FFF9", X"01EC", X"0103", X"008E", X"FFFF", X"FC81", X"FEEB", X"FE48", X"FE40", X"FBA7", X"FC78", X"FFAE", X"01BF", X"FFDF", X"FF8B", X"FB14", X"FF69", X"FF26", X"FEC6", X"FCFD", X"FE24", X"FEA2", X"FCA7", X"FDEA", X"FBEB", X"FC49", X"FBEA", X"FD9F", X"FFF2", X"00C5", X"010D", X"00C6", X"01AA", X"FF08", X"FFBA", X"0016", X"FD25", X"FF4E", X"FE17", X"FD99", X"FF54", X"FFB1", X"0064", X"FC3E", X"01A1", X"FE19", X"FEBB", X"FC82", X"FD2F", X"FCB8", X"FC76", X"FE6A", X"FBFB", X"FC71", X"005F", X"FD96", X"FE5E", X"FDCC", X"FD57", X"FE71", X"FFE3", X"FE03", X"FEFB", X"FF00", X"FF1D", X"FC4E", X"FC7E", X"FD23", X"FD2C", X"FD28", X"FC0C", X"FE09", X"FCCB", X"FDC5", X"FD6D", X"FD47", X"F9ED", X"FB3B", X"FB78", X"FC59", X"FB87", X"FBB9", X"FCD5", X"FDE1", X"FD0B", X"FE1E", X"FE95", X"FE34", X"FEF6", X"021A", X"0306", X"01F1", X"FF1B", X"FB4B", X"FB76", X"FA70", X"FD7E", X"FB98", X"FA18", X"F97C", X"FB98", X"0012", X"FDCE", X"FD6A", X"F6B6", X"FA2A", X"FA52", X"F9D6", X"FA88", X"FD6D", X"FE0C", X"FD5E", X"FD63", X"FE81", X"FEF4", X"FC93", X"00DB", X"04D4", X"043E", X"0222", X"FE97", X"FF00", X"FA9D", X"FB1B", X"FB90", X"F750", X"F8CA", X"F951", X"FB65", X"FFB9", X"FEFF", X"FAE3", X"F890", X"FA1A", X"F9F6", X"FACD", X"FB8E", X"FEA9", X"01A4", X"006A", X"FF63", X"008D", X"FF47", X"FFC4", X"04E5", X"0672", X"075D", X"0427", X"0005", X"FFFB", X"FDEC", X"FF16", X"F915", X"F604", X"F556", X"F6E7", X"F91C", X"FF82", X"FEE8", X"FBCB", X"F978", X"F7FF", X"FAE9", X"FA26", X"FD61", X"01DA", X"0382", X"026A", X"037C", X"01C8", X"0231", X"0518", X"04B4", X"0642", X"0563", X"05A2", X"035A", X"037D", X"00EC", X"FF55", X"FA4C", X"F73E", X"F71F", X"F913", X"FB46", X"010F", X"0079", X"FE27", X"FC59", X"F9DB", X"FBCB", X"FD82", X"FF82", X"01A9", X"0378", X"02CE", X"030B", X"0088", X"02E9", X"0648", X"0643", X"0659", X"0670", X"05A6", X"0641", X"02EF", X"000D", X"FEE6", X"FB33", X"F662", X"F59A", X"F7D8", X"F949", X"FF17", X"FF61", X"FEA5", X"FCF0", X"FC4A", X"000F", X"FDBB", X"FEE8", X"00CB", X"0124", X"01A1", X"017B", X"FEB0", X"02FA", X"050D", X"03ED", X"0474", X"0589", X"055A", X"065B", X"0298", X"FEFE", X"FAD5", X"F851", X"F66B", X"F858", X"F7F5", X"F990", X"FF52", X"FE06", X"008C", X"FE73", X"FF6B", X"FF4E", X"FB5E", X"FB16", X"FE08", X"00F4", X"0043", X"0078", X"0329", X"02E9", X"03FD", X"0385", X"0216", X"054A", X"0417", X"0219", X"FCC5", X"F9DF", X"F8F1", X"F98E", X"F964", X"F4E5", X"F788", X"FBFC", X"FE49", X"005B", X"FED8", X"FE61", X"FBD1", X"FD23", X"F985", X"F935", X"FBE6", X"FECA", X"FF91", X"FF6D", X"00EA", X"0179", X"01C8", X"0489", X"01F2", X"0117", X"029E", X"FD6A", X"FA1A", X"F69A", X"F8F6", X"F8CD", X"F630", X"F882", X"F7F8", X"FA74", X"FE76", X"0074", X"0145", X"FF7D", X"FB07", X"F983", X"F7BA", X"F440", X"F6CD", X"FC10", X"FC66", X"FF72", X"FE3E", X"0167", X"034C", X"02A2", X"004A", X"FCA8", X"FB03", X"F96F", X"F6BB", X"F620", X"FA6B", X"F7F0", X"F846", X"F82F", X"F8C3", X"FCC0", X"FD12", X"FDF2", X"0062", X"FC9D", X"FC3C", X"F9BD", X"F6B3", X"F29C", X"F5F3", X"F90E", X"FB23", X"F8DF", X"FDBE", X"FF90", X"0117", X"016F", X"FD40", X"F914", X"F670", X"F8D6", X"F7AF", X"F71C", X"F7EE", X"F79A", X"F8C0", X"F721", X"F9A2", X"031A", X"00F6", X"0039", X"FDF5", X"FDA9", X"FEB5", X"F995", X"F81C", X"F881", X"F95B", X"F9CC", X"F990", X"FB0B", X"FAB8", X"FC37", X"FE83", X"FE8C", X"FBCD", X"FBDC", X"F854", X"F73B", X"F6DC", X"F611", X"F8C9", X"F903", X"F967", X"F950", X"FC9E", X"0191", X"02C7", X"FF85", X"FD83", X"FBBC", X"FB0C", X"FBC9", X"FBE7", X"FD3C", X"FBFE", X"FC95", X"FBE5", X"FD27", X"FB1E", X"FDFB", X"FC44", X"FB62", X"FBF4", X"FDA6", X"FCB2", X"FB26", X"F99E", X"F71A", X"FA1A", X"FC31", X"FA32", X"FB03", X"FE20", X"00AC", X"005F", X"FFD7", X"00D9", X"FBCD", X"FC9F", X"FE04", X"02D1", X"009D", X"FF72", X"00E0", X"FFE7", X"FF71", X"FD62", X"FB0E", X"FA00", X"FC66", X"FD8F", X"FDE8", X"FEB9", X"FC8B", X"FCDD", X"FCD4", X"FAAD", X"FAA7", X"FE1D", X"FF56", X"00AF", X"FD9E", X"0026", X"0122", X"0106", X"FD9F", X"FE7E", X"0156", X"06ED", X"04C5", X"02D5", X"FFEA", X"024B", X"FFD7", X"FD30", X"FC77", X"FB65", X"FD14", X"FD1D", X"0012", X"02E9", X"01B0", X"0110", X"FDFC", X"FCF1", X"FBCC", X"0053", X"FF7C", X"0062", X"02D8", X"00AF", X"00E3", X"FF01", X"FD4B", X"FD59", X"FE2C", X"06A1", X"03EE", X"021A", X"013C", X"0145", X"0240", X"FFB3", X"FF8A", X"FE6B", X"FDBE", X"001F", X"0230", X"0551", X"0332", X"0124", X"0016", X"FFDB", X"FFAD", X"008E", X"01B0", X"01A0", X"02F2", X"FF8F", X"FEE0", X"002A", X"FDF0", X"FADB", X"FF55", X"04CC", X"00F9", X"0082", X"FE21", X"FD61", X"FDE1", X"FD28", X"FB53", X"FB0E", X"FC9B", X"FB46", X"FD92", X"FEDF", X"0238", X"FFE6", X"FF36", X"02DF", X"026F", X"0343", X"FFFB", X"02AE", X"FFF8", X"000C", X"FF34", X"FFB0", X"00D3", X"0528", X"025D", X"0359", X"FF41", X"FFCE", X"FF90", X"FD3B", X"FC6E", X"FBDC", X"FBCA", X"FBC3", X"FC3D", X"FA56", X"FB11", X"FBE6", X"FDE0", X"FD94", X"FFA7", X"005A", X"006C", X"0332", X"005B", X"00C9", X"FF0D", X"01FA", X"FFC1", X"0077", X"005B", X"FF9E", X"0302", X"051F", X"0505", X"029B", X"0010", X"FFBE", X"00DE", X"FE55", X"FCD7", X"FD30", X"FD0F", X"FE07", X"FD89", X"FE06", X"FD35", X"FCA4", X"FEB9", X"FFD3", X"FDF2", X"035B", X"0293", X"00B8", X"FFB1", X"FF71", X"FFF5", X"FFA9", X"FFD4", X"0008", X"0025", X"FE20", X"FD20", X"FE5B", X"FE6A", X"FCDA", X"FBA1", X"FE04", X"FE9E", X"FAE4", X"FDD0", X"FF6E", X"FA91", X"FAD0", X"FC74", X"FD28", X"FE94", X"FD82", X"FF02", X"006E", X"00EA", X"00B4", X"FF3A", X"00D7"),
--        (X"008C", X"000D", X"FFD8", X"FF7A", X"FF79", X"FF6A", X"00EA", X"003B", X"008D", X"FFF2", X"FF62", X"003F", X"01D9", X"FF82", X"FF67", X"FF92", X"FEEE", X"FF7F", X"0033", X"005C", X"0126", X"0088", X"0102", X"0145", X"FF79", X"FF3B", X"0012", X"00A1", X"FF38", X"0170", X"00F4", X"FFFB", X"00AD", X"0163", X"FE34", X"FD6C", X"0223", X"0157", X"00B1", X"0489", X"0549", X"0355", X"FFD5", X"FF9D", X"FEE6", X"00DB", X"01B7", X"0002", X"0116", X"FED9", X"FF06", X"FEA8", X"006E", X"FF26", X"0031", X"0018", X"007D", X"FF27", X"FF91", X"FF7C", X"00A5", X"0052", X"FF37", X"FDC5", X"0070", X"FEC1", X"FEB7", X"0080", X"0275", X"FF34", X"FFE8", X"FF60", X"008E", X"0546", X"055E", X"0382", X"01A5", X"0038", X"FF88", X"FD14", X"FF73", X"0089", X"000B", X"00C2", X"FF79", X"FF5F", X"0004", X"FD71", X"FFD7", X"0169", X"FF22", X"FF9F", X"0168", X"FFF7", X"038B", X"0254", X"FEC6", X"0022", X"0418", X"034A", X"02EB", X"0598", X"069A", X"0A43", X"07DB", X"07C0", X"0695", X"0248", X"002D", X"FF23", X"FF6E", X"FF05", X"00D0", X"FF2A", X"FE14", X"FC0B", X"FE08", X"0321", X"0363", X"0523", X"0612", X"06C5", X"04E3", X"0108", X"004B", X"00DD", X"03E0", X"04DF", X"08B5", X"082A", X"0483", X"048C", X"08A5", X"08FB", X"0859", X"05A7", X"0239", X"01DC", X"FFDD", X"FFC0", X"00AD", X"FE73", X"FEEA", X"00B9", X"0342", X"0242", X"0548", X"040E", X"061D", X"06A8", X"05B7", X"00D9", X"02C9", X"02D7", X"0475", X"0645", X"08E9", X"06E0", X"0365", X"036F", X"04F1", X"063D", X"090A", X"094A", X"07D2", X"0458", X"01B6", X"00B7", X"FEB2", X"FFCD", X"FFC0", X"FF20", X"0451", X"05BC", X"042A", X"0534", X"04C8", X"037D", X"FF34", X"FEAA", X"FDE0", X"FC5B", X"FCDA", X"FD90", X"FDA6", X"FE51", X"FD71", X"012F", X"0027", X"0161", X"0719", X"0B1D", X"0B2F", X"0642", X"05CE", X"0254", X"009A", X"00BD", X"FEBD", X"0100", X"0712", X"070B", X"044C", X"0574", X"0353", X"019A", X"FD94", X"0090", X"FB42", X"FA5D", X"FA1C", X"F777", X"F900", X"FAD7", X"FAB9", X"FF58", X"FF82", X"00F5", X"0511", X"085D", X"0B1D", X"0A66", X"066A", X"0325", X"04D2", X"FDC3", X"FE94", X"016A", X"03BC", X"0496", X"00A3", X"017B", X"FFB4", X"0113", X"0012", X"FD8C", X"FE3A", X"FB9C", X"FA37", X"F890", X"FD1E", X"FD6B", X"002B", X"012F", X"0339", X"0284", X"03D4", X"05DA", X"09DB", X"0AD8", X"072D", X"008B", X"FDE2", X"FC00", X"0110", X"FFF9", X"045B", X"00DA", X"FDDA", X"FD19", X"FFEC", X"FF76", X"FD7A", X"FCE9", X"FAAA", X"F788", X"F714", X"F79C", X"0017", X"FFDD", X"00C5", X"035F", X"0422", X"04DC", X"0417", X"05D7", X"05F2", X"0A47", X"0132", X"FCEB", X"FE4C", X"FDFC", X"FD0A", X"FEEC", X"01AC", X"FF99", X"FB60", X"FCE5", X"FF9E", X"FD45", X"FCC8", X"FD1F", X"FD1F", X"F97E", X"F6C9", X"FADB", X"FE57", X"0128", X"005A", X"0184", X"002E", X"00B4", X"01BE", X"02ED", X"04DE", X"01F1", X"011F", X"FEEA", X"0001", X"FCA1", X"FB11", X"FDAC", X"FE73", X"FC76", X"FD49", X"FD20", X"FCCB", X"002A", X"FEB6", X"FEBD", X"01BD", X"FE43", X"F6FB", X"FB2A", X"FE42", X"FF83", X"FDAB", X"FEC9", X"FB92", X"FBCA", X"FDF0", X"FE6A", X"0448", X"034F", X"032F", X"FD5D", X"FEC7", X"FF0F", X"FC12", X"FDDC", X"FBAD", X"FBF5", X"FDA0", X"FDA8", X"FDAC", X"FFCE", X"029F", X"054B", X"08B1", X"0640", X"FBF4", X"FD88", X"FFAB", X"FC37", X"FC6C", X"FDDC", X"FDB4", X"FEE0", X"FE1C", X"FE0B", X"04DE", X"00E0", X"FE6B", X"FCAF", X"FF80", X"FF93", X"FC99", X"FCD3", X"FB13", X"FC8E", X"FF5E", X"FF06", X"012E", X"0260", X"05B2", X"094C", X"0A76", X"0560", X"FCC8", X"FFE2", X"002E", X"FFFD", X"FE8B", X"FDCA", X"FDC1", X"FF3A", X"01C7", X"01E1", X"0135", X"0088", X"FFD1", X"FC41", X"018B", X"FFA8", X"FE30", X"FE36", X"FC44", X"005A", X"FF35", X"0127", X"0135", X"03A0", X"042A", X"0827", X"075B", X"027B", X"00FF", X"00EE", X"0115", X"FFA0", X"FD7C", X"FFC7", X"FF1D", X"FF3E", X"FDE8", X"FF0C", X"006A", X"FE8C", X"F9F0", X"FE58", X"00A8", X"FF36", X"0353", X"031D", X"FFC6", X"003D", X"FF55", X"024C", X"029F", X"0200", X"021A", X"046E", X"041B", X"02C4", X"02F6", X"020E", X"FFB6", X"FEB9", X"FDE4", X"FFEA", X"FCDC", X"FE15", X"FE2A", X"FDB7", X"FD94", X"FC57", X"F95B", X"FD5B", X"00CE", X"0122", X"00FF", X"0312", X"0081", X"FFB9", X"FFE9", X"00E5", X"FFBD", X"009E", X"FF5B", X"0239", X"025B", X"0265", X"02E1", X"03DE", X"0029", X"002E", X"FEEF", X"FECA", X"0101", X"00DC", X"FE7E", X"00AB", X"002D", X"FD75", X"FD22", X"FD92", X"FF2E", X"FDB9", X"033B", X"016C", X"0270", X"0259", X"0021", X"007B", X"FEDB", X"FDE9", X"001B", X"022F", X"00ED", X"001D", X"0093", X"01FD", X"0228", X"009D", X"00A5", X"FEFE", X"FF4A", X"FEF2", X"FD67", X"FEF1", X"FDF4", X"F96B", X"FA89", X"FD72", X"FD54", X"00AD", X"012B", X"01A3", X"0262", X"02FF", X"0123", X"0293", X"0198", X"02AA", X"0026", X"00C1", X"034C", X"00B6", X"0099", X"FFCB", X"0073", X"FFA4", X"FF69", X"FE36", X"FE0B", X"FDB2", X"FD7F", X"006B", X"FC96", X"F9DE", X"FAB2", X"FB7C", X"FF30", X"FFB3", X"FEFB", X"FF9F", X"013A", X"037E", X"0237", X"03F5", X"02E5", X"0176", X"03EF", X"03F5", X"00E7", X"FCFB", X"FF3B", X"0070", X"0103", X"0134", X"0273", X"FF10", X"FED2", X"01C4", X"0114", X"FF73", X"FCA8", X"F7F0", X"FBDD", X"FDE4", X"00CB", X"0227", X"043D", X"02AE", X"0253", X"065D", X"07F1", X"088A", X"06AF", X"0528", X"020B", X"02A8", X"013B", X"FF46", X"FEA9", X"00C9", X"00D0", X"02D1", X"04B2", X"0109", X"02AD", X"00BB", X"0177", X"FEE9", X"F902", X"F8D7", X"FE4A", X"FFD4", X"0146", X"0081", X"0400", X"0559", X"034E", X"07F2", X"08A9", X"08D8", X"060D", X"01D1", X"00F4", X"01EF", X"0047", X"FFDF", X"0352", X"0176", X"01BC", X"030E", X"0320", X"003E", X"00AD", X"014D", X"0219", X"FFDC", X"FBEA", X"FCF0", X"025B", X"FF70", X"FF27", X"FFB9", X"032D", X"0461", X"0204", X"04C1", X"0895", X"0807", X"03A0", X"007B", X"00CF", X"02B2", X"0275", X"03D3", X"0156", X"00DF", X"026A", X"02B0", X"0341", X"055B", X"011F", X"02AE", X"02F6", X"FE51", X"FBF8", X"FC51", X"01B9", X"FF58", X"0037", X"00E8", X"03C8", X"0432", X"0067", X"FFE8", X"0228", X"026F", X"021A", X"01BF", X"035E", X"0343", X"0374", X"037E", X"036B", X"030B", X"03C5", X"031F", X"0538", X"0396", X"0360", X"00D1", X"0019", X"FE9B", X"FC5B", X"FED2", X"FE9A", X"FF93", X"FE83", X"0076", X"FEE9", X"0130", X"FBD2", X"F7D3", X"FA95", X"FD92", X"FE6D", X"006F", X"0103", X"028D", X"01D5", X"03DF", X"036A", X"022D", X"02F9", X"FFF8", X"FFE0", X"00AD", X"FD8F", X"FD0D", X"FEFB", X"FFE4", X"FF53", X"023B", X"00AC", X"0058", X"FF77", X"FE93", X"FF1B", X"FF25", X"F9C2", X"F686", X"F8BD", X"FA12", X"F86E", X"FB66", X"FD32", X"FCBD", X"FAE7", X"FD22", X"FD56", X"FFC7", X"FE0D", X"FB9D", X"FC4E", X"FBCF", X"FB9A", X"FB3E", X"FE05", X"011D", X"0012", X"FEDD", X"0234", X"FF90", X"00E6", X"00B6", X"0081", X"FE59", X"FC5E", X"FA7A", X"F71E", X"F798", X"F672", X"F4D7", X"F69E", X"F7E7", X"F870", X"F5F5", X"F2BB", X"F784", X"F992", X"F921", X"F91F", X"F934", X"FB9A", X"FB61", X"FB2E", X"013D", X"FEB1", X"FFD7", X"00A8", X"0141", X"0017", X"FFA8", X"FFEC", X"FF95", X"FFAE", X"FF72", X"FC91", X"FCEB", X"FD1A", X"FB12", X"FC93", X"FE48", X"FDF7", X"FCB0", X"F682", X"FAD9", X"FB30", X"FBC0", X"FC13", X"FC33", X"FFB8", X"FBFD", X"FDA7", X"FE66", X"FEEA", X"015D", X"0044", X"0130"),
--        (X"FF4B", X"FF0D", X"FF51", X"FFDE", X"FF9B", X"FF98", X"00D9", X"0187", X"FF30", X"FF58", X"00B0", X"006A", X"FEF6", X"FDA3", X"FF8F", X"FF10", X"FF42", X"FFCF", X"0069", X"004D", X"FFB9", X"0050", X"FE3E", X"0096", X"001F", X"0043", X"00B2", X"FFAB", X"FF92", X"0022", X"0083", X"FF83", X"0108", X"FEC6", X"FC28", X"FB3E", X"FC16", X"FB6D", X"FA81", X"FA8A", X"F8DB", X"F6B4", X"F9EC", X"FD17", X"FF87", X"FD2F", X"FB5D", X"FC5C", X"FD21", X"FF24", X"FF23", X"FE30", X"FF55", X"00DC", X"FF81", X"0110", X"0008", X"FF5F", X"0061", X"FF01", X"FE0F", X"FCF5", X"F9EE", X"FA74", X"F92A", X"FB9C", X"F9E7", X"FB40", X"FCF2", X"FD26", X"FA45", X"FCE9", X"FB96", X"FC56", X"FE99", X"FAB8", X"FC0E", X"FBF7", X"FB10", X"FEBA", X"012A", X"0040", X"005D", X"FFC3", X"FE1B", X"FFE4", X"0074", X"FD8B", X"FC28", X"01D0", X"0075", X"00CF", X"FF12", X"FFE4", X"FC90", X"FEEF", X"008E", X"FD39", X"FD4A", X"FD97", X"FE20", X"FDCA", X"FF2F", X"FCD2", X"FAF9", X"F98E", X"FB70", X"FAB2", X"FD2F", X"FF0D", X"FF18", X"FFE9", X"FF90", X"FFDE", X"FF55", X"00DB", X"01ED", X"0444", X"025F", X"00EF", X"0316", X"0279", X"FFF4", X"FFFB", X"FF03", X"00CB", X"0118", X"FFDA", X"FF8F", X"FEE7", X"FED8", X"FEF1", X"FE22", X"FC1C", X"F9F8", X"F73A", X"FB57", X"FCC5", X"011C", X"FFA6", X"FECF", X"FF35", X"007B", X"02FE", X"046D", X"04A2", X"020C", X"001C", X"FD97", X"FF25", X"FE40", X"FEB9", X"00AF", X"01CA", X"015C", X"0540", X"03E8", X"0018", X"FE84", X"FE1C", X"FF24", X"FDD5", X"F975", X"FAB4", X"FB42", X"FE73", X"0127", X"FF5E", X"006C", X"FEAE", X"FCAC", X"FFF1", X"01B4", X"0076", X"FF5B", X"FFC8", X"FE6D", X"FDDA", X"0001", X"0096", X"FF41", X"01C8", X"05AF", X"07D8", X"0646", X"029B", X"FEEE", X"FDB0", X"FDAE", X"FCC3", X"FA2B", X"FB2C", X"F8A2", X"FCD8", X"FEFB", X"FFE1", X"FF3B", X"0145", X"FD88", X"FE6C", X"0320", X"FFE0", X"FD90", X"FCB2", X"FCCB", X"FC71", X"FDC5", X"FC31", X"005D", X"02A8", X"056E", X"0902", X"0574", X"FEE4", X"FDDC", X"FCBC", X"FEE7", X"FFA4", X"FB4E", X"FD40", X"FB13", X"FB22", X"FF96", X"002F", X"FD9D", X"FAE9", X"FB29", X"FC90", X"00C7", X"FD37", X"FD54", X"FE35", X"FCB1", X"FD4C", X"FBCE", X"FA27", X"FBD0", X"00AF", X"0724", X"07C7", X"04E9", X"FFF9", X"FE7A", X"FF01", X"FDD1", X"FE67", X"FFF1", X"FB77", X"F91D", X"FCED", X"FF4D", X"028A", X"FF5C", X"FB48", X"FCBB", X"FC6F", X"FF8C", X"FF19", X"FFE7", X"003F", X"FDCA", X"FC5C", X"FACC", X"F70F", X"F903", X"008B", X"08D3", X"09C8", X"0517", X"02B5", X"000A", X"018D", X"01BD", X"0157", X"0369", X"FF9D", X"F956", X"F708", X"FDD8", X"FFCE", X"FEA3", X"FBB6", X"FA1B", X"FE82", X"0015", X"0052", X"0222", X"00C9", X"FE08", X"FB3B", X"F94D", X"F6CB", X"F9B2", X"01C1", X"0A91", X"0981", X"0657", X"0195", X"012A", X"028A", X"0273", X"0234", X"03F6", X"02E4", X"FD74", X"F7BC", X"FC25", X"0126", X"FE62", X"FB9C", X"F7E0", X"FEE6", X"FF3C", X"0295", X"0016", X"FF23", X"FF0F", X"FBCF", X"F9E9", X"F68A", X"FAD4", X"0428", X"0CF3", X"08BE", X"021D", X"FFE1", X"0221", X"030E", X"0422", X"05AA", X"0570", X"0265", X"FFC3", X"FE5A", X"002D", X"0086", X"FE93", X"F92C", X"F6E7", X"FBC2", X"008C", X"FE46", X"FCF0", X"FC9C", X"FD72", X"FD02", X"FA53", X"F7F9", X"FD02", X"07FA", X"0A5D", X"040E", X"016B", X"FFAB", X"009B", X"02CF", X"04E0", X"04F3", X"03AF", X"004B", X"FE3B", X"00BE", X"01F1", X"01CD", X"0041", X"FD22", X"F9DD", X"FE5D", X"002B", X"FD19", X"FC0D", X"FDCA", X"FD5A", X"FBB9", X"FAD8", X"FB40", X"03EA", X"087C", X"08ED", X"0443", X"01C0", X"012F", X"01F3", X"034C", X"015D", X"00CF", X"FD9A", X"FB53", X"FBEC", X"020E", X"072A", X"0424", X"FDF7", X"FE1A", X"F8DB", X"FDEF", X"FEC2", X"FBC2", X"FBFE", X"FD16", X"FD22", X"FC86", X"FDCD", X"FE11", X"05A1", X"094E", X"0822", X"028C", X"0022", X"026E", X"00AE", X"016F", X"0178", X"FEC0", X"FDD4", X"F998", X"FAC0", X"041A", X"07B7", X"0445", X"FD9B", X"0012", X"FA47", X"FFAF", X"00CE", X"FFE2", X"FED5", X"FD67", X"FE21", X"FDF8", X"FF8E", X"02B6", X"0533", X"0895", X"06C2", X"0273", X"01C5", X"00C0", X"0257", X"0021", X"FFB0", X"FD51", X"FC18", X"F981", X"FCA0", X"052B", X"05BB", X"0230", X"0053", X"FFC9", X"FFBD", X"00E0", X"0222", X"0040", X"FE98", X"FF64", X"FDAE", X"008F", X"004D", X"0458", X"070E", X"0925", X"03C4", X"003E", X"0294", X"02EB", X"FF77", X"FB67", X"FE58", X"FD6D", X"FD4B", X"FE33", X"FFB9", X"059D", X"07E3", X"0347", X"FFD0", X"02BB", X"0067", X"03BA", X"023B", X"009A", X"FF1A", X"FF74", X"FFB5", X"009A", X"00C7", X"042C", X"0848", X"06B0", X"0126", X"0260", X"01F3", X"00A2", X"FD35", X"FD98", X"FE07", X"FD88", X"FEA1", X"FD96", X"FFD9", X"0796", X"05F9", X"01D8", X"FE88", X"FFEF", X"FC8C", X"00E6", X"0003", X"0237", X"0074", X"00FC", X"0019", X"002F", X"0204", X"05F2", X"06CF", X"0406", X"009B", X"02CE", X"033D", X"013B", X"FFAC", X"FE61", X"FD75", X"FF6B", X"0040", X"0205", X"FFE0", X"02CE", X"02B8", X"03A7", X"FF46", X"FAF5", X"FDEE", X"FF5D", X"FF27", X"01D9", X"0001", X"04A1", X"0143", X"0251", X"06F2", X"0510", X"0324", X"023C", X"0096", X"0280", X"025F", X"FEED", X"FEFD", X"0057", X"FFC2", X"FEFB", X"014D", X"0245", X"FFE6", X"03BE", X"05AE", X"02B2", X"0021", X"FED1", X"0084", X"FF3E", X"00BC", X"01A0", X"035F", X"0339", X"0220", X"0374", X"02AF", X"0087", X"FDF0", X"FC80", X"FE89", X"005F", X"FFB0", X"FF43", X"FE33", X"0002", X"FF7B", X"001E", X"0025", X"00D2", X"01DA", X"023F", X"0064", X"0155", X"FFCB", X"0071", X"01FF", X"016D", X"0010", X"01A4", X"03D7", X"044A", X"02AA", X"02E2", X"0104", X"FE91", X"FDC1", X"FCD0", X"FE34", X"FCD4", X"0041", X"FE74", X"FF25", X"001B", X"FF03", X"FDE6", X"FF0E", X"0131", X"03CB", X"0039", X"FDDB", X"00D5", X"007B", X"0095", X"0469", X"0262", X"01CB", X"0235", X"03E6", X"049D", X"0227", X"0265", X"0095", X"FF3D", X"FFC5", X"FE7C", X"FD9C", X"FC50", X"FCE9", X"FEC9", X"FE32", X"FD0E", X"FDCD", X"FD98", X"0024", X"00C8", X"01D0", X"00FC", X"FD81", X"FFC8", X"FFAA", X"FF78", X"0270", X"01A8", X"0207", X"005D", X"01FB", X"023C", X"027A", X"0079", X"FF38", X"FFD3", X"FF33", X"FD5A", X"FCA9", X"FD71", X"FCEA", X"FE30", X"010E", X"FF5C", X"00ED", X"0162", X"0201", X"020A", X"01D7", X"FF2D", X"FD6C", X"0008", X"FEB8", X"FEF3", X"0113", X"000B", X"FF78", X"000B", X"0257", X"019B", X"FF89", X"FEE0", X"FE6E", X"FE0E", X"FD45", X"0009", X"FE26", X"FE33", X"FFD1", X"FEE1", X"FF21", X"0199", X"0209", X"0251", X"03C2", X"0449", X"FFB1", X"FF24", X"FF9C", X"00C1", X"00D3", X"0050", X"022C", X"FD95", X"FFAF", X"0127", X"0090", X"FE6B", X"FCDA", X"FBBF", X"FE5A", X"FD05", X"FDBB", X"FDFA", X"FF9A", X"FD05", X"FF32", X"FF67", X"FF52", X"00E1", X"026D", X"0300", X"FDEF", X"0073", X"FD48", X"0213", X"0059", X"00BB", X"000E", X"00F3", X"004B", X"000D", X"0164", X"00C8", X"01DF", X"0012", X"FE05", X"FE43", X"FF3D", X"0041", X"FF4D", X"FFA4", X"0217", X"FE30", X"01AF", X"011E", X"009C", X"FE23", X"009A", X"02C0", X"0188", X"032D", X"0224", X"FEA2", X"FEF1", X"FEDB", X"0006", X"FEF6", X"002E", X"FFB3", X"FD32", X"FE85", X"00BF", X"FFAA", X"FE4E", X"FC1B", X"FC9F", X"FDCF", X"FDB1", X"FA37", X"005F", X"001D", X"FEDF", X"FD58", X"FDBF", X"FC86", X"FEEB", X"FE16", X"FF0F", X"FBAB", X"FF10", X"FF55", X"007C", X"0059"),
--        (X"FF17", X"FEB2", X"00A3", X"FF75", X"0031", X"00BF", X"008F", X"0105", X"FEB6", X"FF0A", X"017C", X"0012", X"FF77", X"0076", X"0186", X"0222", X"00E8", X"FFA8", X"FF54", X"FFD4", X"FEDD", X"FFC4", X"0165", X"0042", X"0040", X"0163", X"0075", X"00EA", X"FE0F", X"FFAF", X"FE59", X"0156", X"FF6C", X"FF13", X"FDE5", X"0006", X"FF84", X"FEF5", X"FE83", X"0000", X"0050", X"FE60", X"FCE2", X"FBF6", X"FF2B", X"0001", X"FDFF", X"FEE9", X"FF3B", X"FFC8", X"FEA5", X"0060", X"004A", X"FF23", X"0121", X"00D3", X"00A8", X"00E5", X"FEFB", X"01DC", X"0006", X"FF3E", X"FD89", X"FD95", X"FD4E", X"FE5D", X"FBE5", X"FE93", X"FB29", X"FA59", X"FB4D", X"FAFA", X"FCEE", X"FEFC", X"FECF", X"FDF0", X"FF03", X"FF3C", X"00A4", X"0059", X"0272", X"03B5", X"005C", X"0013", X"FEFC", X"0067", X"FEE2", X"FEAF", X"FED3", X"FCD8", X"FE2C", X"FF0E", X"FEE3", X"FE5A", X"0236", X"024F", X"02B2", X"00D7", X"0221", X"0223", X"0198", X"00D1", X"FFC6", X"00EC", X"035F", X"0309", X"0218", X"0154", X"013D", X"01EE", X"00ED", X"0091", X"0052", X"FFBC", X"FF65", X"0157", X"FE49", X"FE3B", X"FEEC", X"FE5D", X"FE99", X"02A0", X"0260", X"052A", X"045E", X"01D9", X"046F", X"04C0", X"0212", X"FEE6", X"FE45", X"FDF7", X"FEA3", X"FF4D", X"FBE9", X"FD71", X"016A", X"046D", X"0309", X"FE12", X"001F", X"01FD", X"FFE4", X"02CA", X"FEB0", X"0105", X"00A7", X"02C6", X"0453", X"05EB", X"0511", X"06B3", X"0746", X"05E9", X"0574", X"038E", X"0416", X"02D6", X"008A", X"FEAC", X"FE52", X"FE5B", X"FD95", X"FC60", X"FBDA", X"07B8", X"028A", X"FD56", X"FED8", X"012C", X"023C", X"0322", X"00EE", X"03F4", X"054A", X"065F", X"08DE", X"084F", X"0693", X"087F", X"065F", X"0699", X"0471", X"0331", X"033B", X"0246", X"0149", X"0009", X"0045", X"01A8", X"FFD3", X"FDF1", X"FFB2", X"0302", X"0375", X"FF7A", X"018D", X"031E", X"0394", X"052E", X"03F9", X"0618", X"0803", X"08E8", X"0979", X"0883", X"076C", X"03C8", X"0499", X"01EB", X"00CC", X"0113", X"021C", X"01C9", X"0299", X"0175", X"00D5", X"027B", X"01BB", X"0273", X"02E7", X"057D", X"0181", X"0122", X"00F6", X"05AC", X"0156", X"0718", X"0632", X"07CF", X"0954", X"0A6B", X"08FF", X"07FF", X"0456", X"04C1", X"02D7", X"01DE", X"FFC6", X"0421", X"031F", X"02E6", X"0353", X"024C", X"02F5", X"01B6", X"048F", X"0681", X"05EA", X"0484", X"072A", X"052D", X"01AD", X"02AD", X"03A5", X"0951", X"0600", X"080E", X"0828", X"0673", X"0491", X"037F", X"0202", X"01B4", X"02FF", X"0380", X"059A", X"0332", X"045C", X"061C", X"0388", X"0389", X"025D", X"0485", X"0438", X"05AD", X"07E5", X"0B56", X"097F", X"038B", X"003C", X"00A8", X"050D", X"0581", X"0719", X"0612", X"04E0", X"0207", X"00D1", X"0189", X"007E", X"0279", X"0173", X"04CC", X"04C9", X"0199", X"0433", X"044D", X"048E", X"0205", X"0206", X"027B", X"04B2", X"0426", X"0408", X"0762", X"07AF", X"017F", X"00E4", X"032D", X"0785", X"0518", X"03A4", X"0151", X"0176", X"003F", X"FF18", X"FF1F", X"FEAE", X"0062", X"0060", X"03AC", X"FC95", X"FBE5", X"FF42", X"0011", X"0088", X"FF49", X"FE77", X"FEEA", X"FD50", X"FE08", X"FFA9", X"051A", X"039A", X"FDE8", X"00D6", X"03B5", X"0474", X"034B", X"FED6", X"FC54", X"F808", X"FB38", X"FC84", X"FBC6", X"FDE7", X"FDF3", X"FDF8", X"FA70", X"F964", X"FA84", X"FF56", X"FF5C", X"FD45", X"FD21", X"FDDC", X"FBE9", X"FAE9", X"F95B", X"FD9F", X"0178", X"039D", X"FE74", X"FFDB", X"01F1", X"04E8", X"FF53", X"F9D3", X"F7F3", X"F55D", X"F885", X"FAF4", X"FC13", X"FBA6", X"FB2B", X"F9DC", X"F814", X"F861", X"FA73", X"FC7A", X"FDA8", X"FD84", X"FD80", X"FC25", X"FBE6", X"FB3C", X"F9BF", X"FD49", X"FF13", X"03C9", X"0367", X"0267", X"010D", X"0307", X"FE13", X"FB17", X"F7A6", X"F30D", X"F845", X"F979", X"FB75", X"FBC6", X"FDDE", X"FC52", X"F9CB", X"FAF3", X"FA5D", X"FD4A", X"FE6E", X"FFF8", X"FE74", X"FF74", X"FCD9", X"FA59", X"FD15", X"007D", X"0040", X"060E", X"0339", X"00F6", X"FF10", X"03B9", X"0111", X"FF47", X"F969", X"F63D", X"F609", X"F819", X"FC89", X"FCC2", X"FCD6", X"FDA1", X"FD29", X"FAC8", X"FBCA", X"FC64", X"FEF6", X"0239", X"0161", X"FFCB", X"FFED", X"FF16", X"00A1", X"039D", X"01DD", X"04CF", X"03B5", X"01D9", X"FF8D", X"0256", X"02FD", X"02D4", X"FC76", X"F769", X"F7F3", X"F9CD", X"FD6B", X"FCAC", X"FD05", X"FEE3", X"FD07", X"FA55", X"FBEA", X"FC75", X"00E5", X"0236", X"01AA", X"0151", X"012E", X"01BB", X"02B6", X"02EC", X"0388", X"036A", X"04DA", X"001B", X"FFEA", X"011D", X"0378", X"0605", X"009F", X"FC52", X"F6BD", X"F90A", X"FB2C", X"FA7C", X"FC3C", X"FC55", X"FAE5", X"F978", X"FA8E", X"FF50", X"00F2", X"0285", X"012E", X"00E6", X"0197", X"03E8", X"039C", X"045C", X"0459", X"02E8", X"036C", X"00E7", X"FEBF", X"0151", X"0204", X"0498", X"056B", X"0063", X"FBEA", X"FA17", X"FAFD", X"F960", X"FB15", X"FB00", X"FB1F", X"FB18", X"FCC0", X"FF68", X"02E6", X"FFB8", X"00FC", X"015C", X"01B4", X"02B5", X"0501", X"050A", X"01DF", X"0132", X"FFA0", X"FFFD", X"038A", X"01E5", X"009E", X"0643", X"068A", X"044D", X"0184", X"FFB0", X"FE31", X"FE43", X"FD01", X"FEC7", X"FD15", X"FD0C", X"FFCF", X"FEE4", X"0013", X"0012", X"FF0B", X"0096", X"02CB", X"028B", X"0477", X"02F9", X"00BE", X"009A", X"FEAB", X"00D7", X"0054", X"0309", X"023E", X"0763", X"0855", X"070D", X"061C", X"0225", X"01A9", X"015A", X"008E", X"0127", X"0034", X"0007", X"0103", X"FE12", X"FED5", X"FD45", X"FF25", X"FF28", X"024B", X"0446", X"03E2", X"FFF7", X"0135", X"FFDC", X"FDCA", X"FFC8", X"00B3", X"0297", X"056F", X"07A1", X"06B2", X"08E1", X"075A", X"0619", X"04EC", X"0144", X"02F4", X"0229", X"010C", X"FEBF", X"FFB6", X"FF1C", X"0058", X"FE56", X"FDBA", X"FD89", X"017E", X"043F", X"03DF", X"006F", X"0587", X"00FB", X"008A", X"FE9B", X"00C0", X"01E1", X"00F1", X"0387", X"01E7", X"076D", X"097A", X"07A8", X"051A", X"044A", X"043B", X"04F3", X"04C8", X"0133", X"0178", X"FFD2", X"FE01", X"FDCA", X"FCCC", X"FE42", X"0028", X"025C", X"FF8F", X"008A", X"02E3", X"FE7C", X"0021", X"FFF7", X"005E", X"0169", X"04AE", X"0262", X"FCCB", X"00AA", X"044D", X"02AF", X"045D", X"0709", X"07A9", X"0425", X"0391", X"05ED", X"03EB", X"01FF", X"0023", X"FEBE", X"FCC2", X"FBAD", X"FD2F", X"FE57", X"FDC3", X"FFEE", X"00CF", X"FDBC", X"FE95", X"FF5F", X"FF9E", X"0028", X"0647", X"030B", X"FF6D", X"FF88", X"0142", X"026B", X"01BC", X"0239", X"0419", X"06FE", X"082C", X"0740", X"05CC", X"0478", X"020D", X"FFD4", X"FF19", X"FA64", X"FBB3", X"FD23", X"FB55", X"013A", X"FE15", X"FE96", X"FF9C", X"0090", X"FE54", X"FCF9", X"0436", X"0316", X"00D5", X"013C", X"00FC", X"FF73", X"0239", X"023A", X"0379", X"0375", X"01EE", X"02B5", X"0501", X"04A4", X"0362", X"03F1", X"007C", X"FBE2", X"F938", X"FED4", X"FE87", X"0274", X"FFE1", X"00CC", X"FFAE", X"0034", X"FFB3", X"FFF1", X"FDDE", X"FB8C", X"FE9C", X"FF45", X"FE0C", X"0075", X"0119", X"FEF5", X"FFF8", X"FDF1", X"00D7", X"FE87", X"0276", X"0379", X"03C8", X"0549", X"0505", X"0076", X"FED5", X"00FB", X"FFB5", X"007B", X"FEA1", X"FF70", X"FFF1", X"FFD9", X"0083", X"FFD2", X"00C4", X"0124", X"0240", X"01FA", X"0155", X"03D7", X"0236", X"041E", X"0169", X"0172", X"0716", X"031A", X"0086", X"0146", X"047C", X"03E8", X"0541", X"02D3", X"028F", X"01D9", X"03C0", X"FF3D", X"003D", X"FFDD", X"009D"),
--        (X"FF88", X"FF3F", X"FFB9", X"0119", X"FF42", X"00AD", X"FFFE", X"FE19", X"0059", X"00A8", X"FFF0", X"0098", X"0007", X"FF56", X"0044", X"0053", X"0125", X"FFCF", X"0009", X"002E", X"00D3", X"0062", X"FFAA", X"FFC3", X"0019", X"0051", X"020F", X"0055", X"0120", X"FFD7", X"FEE3", X"0043", X"001F", X"FF85", X"012E", X"FF36", X"011B", X"012A", X"0159", X"0170", X"011C", X"00D8", X"FFE2", X"FD99", X"00F6", X"0023", X"00D6", X"036A", X"019F", X"01CF", X"FFE3", X"0181", X"0069", X"006A", X"0035", X"FF89", X"FFEC", X"FE60", X"FFD4", X"0032", X"FEDE", X"0097", X"00BB", X"00BD", X"038D", X"0672", X"0627", X"05B3", X"0618", X"02C8", X"05D1", X"01E0", X"0281", X"01BB", X"019C", X"FF9D", X"0191", X"00FD", X"0134", X"00C9", X"0356", X"03B1", X"000D", X"0096", X"0026", X"0048", X"FC2A", X"014F", X"0094", X"FD4A", X"004A", X"FF0D", X"005B", X"05B2", X"0399", X"025B", X"00D2", X"02C1", X"0233", X"00C6", X"FFBB", X"00C6", X"FF90", X"01F3", X"FEAA", X"FFDA", X"00A1", X"005F", X"0103", X"FE28", X"FF67", X"FF98", X"FF79", X"FF0F", X"FCC3", X"FDB3", X"FF2C", X"FD35", X"FE95", X"FEB8", X"FF5E", X"01DF", X"0093", X"FDF1", X"FEFC", X"00C6", X"FDAE", X"FDBE", X"FEE9", X"0143", X"FC3B", X"FDA2", X"007E", X"0010", X"00A0", X"0180", X"FF5B", X"FD88", X"FD91", X"00AC", X"00C8", X"FEFF", X"FE99", X"FF75", X"FDDF", X"FCEC", X"FE0A", X"002F", X"FFE4", X"0122", X"0150", X"FDCF", X"FF45", X"FD8A", X"0040", X"0003", X"0102", X"FF88", X"0131", X"FF78", X"FFB8", X"FF08", X"FF5B", X"0214", X"FED3", X"FDD3", X"FDC3", X"011C", X"00CE", X"FF35", X"FDFF", X"0049", X"FDF1", X"FD38", X"FE68", X"0285", X"0087", X"00B1", X"FDF6", X"FEF6", X"FEFE", X"FFA1", X"00FA", X"021E", X"0183", X"013E", X"006E", X"FF67", X"0018", X"030A", X"00CB", X"FEB5", X"FD39", X"FB3D", X"F8D2", X"FE5F", X"0034", X"FFFB", X"0423", X"01D0", X"FEEA", X"FD67", X"0043", X"0031", X"FE62", X"FFAA", X"0076", X"01D2", X"FFB6", X"0111", X"00E3", X"00CC", X"0247", X"012E", X"01FB", X"FFFE", X"0031", X"00C6", X"01F0", X"FF9D", X"FE1F", X"F7EC", X"F9C4", X"FF52", X"0191", X"0576", X"0230", X"0136", X"FED1", X"FE21", X"FD8A", X"00FE", X"0048", X"0018", X"00C3", X"011E", X"00FF", X"0111", X"029D", X"020F", X"0251", X"027D", X"0051", X"FFC7", X"00DA", X"FE95", X"0080", X"FEEB", X"FBC4", X"F730", X"FAF0", X"FCDF", X"0270", X"050E", X"00BC", X"00DE", X"FF58", X"FFEA", X"FEE8", X"FEAE", X"FDD6", X"FE7B", X"FFF3", X"FFC0", X"FFE8", X"0026", X"FFA7", X"00AB", X"045C", X"021B", X"021B", X"0020", X"FFD3", X"FEFE", X"FF48", X"FDB4", X"FA8C", X"F56B", X"F89C", X"0028", X"025F", X"0346", X"04BB", X"01DD", X"FF57", X"0381", X"00F5", X"0034", X"FEB8", X"FE00", X"FE7A", X"FD8B", X"FC92", X"FD59", X"FB1D", X"FCE0", X"0335", X"018D", X"02D8", X"00FA", X"FF64", X"00BD", X"0187", X"FD69", X"F924", X"F64A", X"F764", X"FC00", X"0204", X"047B", X"06BE", X"036D", X"02DB", X"0324", X"02EE", X"FFB3", X"FED4", X"FD52", X"FF0E", X"FE72", X"FA69", X"FBB7", X"F92D", X"FA39", X"FE21", X"FFAB", X"00A6", X"0042", X"00E6", X"017A", X"0338", X"010F", X"F9D6", X"F560", X"F950", X"FE98", X"006E", X"03C6", X"098E", X"0884", X"043E", X"0487", X"0121", X"0041", X"FEF3", X"FC94", X"FBD8", X"FC93", X"FC8A", X"FA46", X"F747", X"FA20", X"FD54", X"FDAA", X"FE4D", X"FEDB", X"FFE3", X"031C", X"0689", X"05D0", X"0990", X"02D8", X"0116", X"0298", X"FEFD", X"03BE", X"080E", X"0980", X"0876", X"0791", X"06CD", X"02C6", X"0027", X"FB3C", X"FD82", X"FBFC", X"FA9D", X"F95F", X"F94F", X"FA12", X"FA73", X"FDC7", X"FE91", X"FF69", X"FF1E", X"0439", X"0562", X"064B", X"0A8F", X"0A63", X"051C", X"02C1", X"FE98", X"FF4B", X"0484", X"05A1", X"0827", X"0945", X"0A24", X"0864", X"03D3", X"0171", X"FF51", X"FC95", X"FB28", X"FA7B", X"F9E3", X"FA40", X"FB6C", X"FE79", X"0170", X"034E", X"0353", X"025A", X"02A2", X"03EA", X"0490", X"0670", X"0745", X"0370", X"0121", X"FE36", X"FD81", X"0313", X"0647", X"09EA", X"0ADC", X"0ADA", X"0898", X"0663", X"044B", X"000A", X"FA29", X"F9F4", X"F9B6", X"FDE7", X"007B", X"040F", X"02AD", X"0431", X"0382", X"0205", X"FEA1", X"FFA5", X"FFA8", X"03E7", X"0729", X"039C", X"015F", X"FE41", X"FE77", X"FF16", X"0161", X"02B7", X"05E4", X"0851", X"0868", X"0759", X"0774", X"044C", X"0113", X"FEA8", X"FF68", X"006F", X"021C", X"0494", X"02CF", X"03E8", X"02CD", X"0072", X"FF09", X"FC50", X"001C", X"0A70", X"0723", X"0222", X"0113", X"FD5B", X"0099", X"FC42", X"FD63", X"FFB2", X"FEE3", X"01E7", X"0635", X"076C", X"0BAF", X"0AFC", X"0519", X"044B", X"0225", X"00FB", X"0025", X"0136", X"0197", X"00CC", X"003C", X"FF29", X"FE4F", X"FB85", X"00D3", X"0C70", X"0798", X"050B", X"02C7", X"FE83", X"FFD6", X"FE7A", X"FE2F", X"FE88", X"FCF6", X"FFEB", X"0110", X"048E", X"087A", X"082D", X"086B", X"04F5", X"FFDD", X"FF87", X"FFF2", X"0018", X"FFEF", X"01C9", X"FF11", X"FE7C", X"FDD1", X"FFF8", X"040A", X"09BA", X"03BC", X"0190", X"006A", X"01E9", X"0167", X"FEEC", X"FDDE", X"FC53", X"FC8D", X"FED2", X"FF31", X"0184", X"020C", X"0601", X"05A4", X"037E", X"02A0", X"FE50", X"FE3C", X"00A3", X"FEC6", X"FDC8", X"FE89", X"FE28", X"FE46", X"0025", X"03CB", X"0591", X"02D0", X"0211", X"0136", X"0033", X"0151", X"00B1", X"FF80", X"FE97", X"FD1D", X"FEAE", X"FE00", X"FDE3", X"0006", X"01C5", X"05C8", X"02B6", X"0217", X"012D", X"0036", X"FE95", X"FECF", X"FEA4", X"FE30", X"FF45", X"FDA4", X"FF79", X"05C8", X"04F6", X"013F", X"FE61", X"FE96", X"FEC7", X"00F4", X"FF69", X"FBB9", X"FF11", X"FD14", X"FD66", X"FE92", X"FE7A", X"FEFD", X"004C", X"018E", X"0232", X"0101", X"00CC", X"003C", X"FF24", X"FF2F", X"FF08", X"00C0", X"003D", X"0254", X"082C", X"060E", X"075B", X"03E3", X"006F", X"FF09", X"00D9", X"0004", X"FCF1", X"FE56", X"FF18", X"FF6E", X"FF5A", X"004B", X"FF96", X"009E", X"FE90", X"0000", X"0052", X"FF80", X"002B", X"0013", X"FE10", X"00DF", X"0166", X"00E2", X"01C7", X"04FA", X"0695", X"07DB", X"04BE", X"FF5B", X"0118", X"FF25", X"FF59", X"FC90", X"FA61", X"FA17", X"FF42", X"0104", X"0171", X"0100", X"FFF7", X"FEBE", X"006F", X"0109", X"01E8", X"0099", X"00C4", X"000F", X"FF04", X"00C9", X"01FD", X"002F", X"069E", X"0729", X"060E", X"03D5", X"0543", X"FF8B", X"FFDA", X"0003", X"0112", X"FD9E", X"FA2D", X"FE25", X"027E", X"0015", X"FEA4", X"FF00", X"FE17", X"FD60", X"FE3D", X"FF3D", X"FF0F", X"00F1", X"0066", X"FCAD", X"FCBB", X"FE2E", X"FE48", X"FE92", X"0372", X"03CF", X"0194", X"045D", X"04B5", X"00D1", X"0082", X"FF87", X"FE96", X"FE89", X"0129", X"02E5", X"013B", X"FFC7", X"FFEC", X"FE6D", X"FC3E", X"FC51", X"FD74", X"FD93", X"FE13", X"FF65", X"005F", X"FCFB", X"F9A8", X"FB89", X"FAEA", X"FC4E", X"FE7C", X"FC4E", X"FC24", X"FCA6", X"0168", X"0251", X"0035", X"FF0B", X"FFC0", X"FEF4", X"001C", X"FFAE", X"00FC", X"02A0", X"0322", X"023B", X"022B", X"0172", X"0257", X"04B5", X"0707", X"07A8", X"064F", X"0370", X"031A", X"023C", X"0385", X"00E6", X"FFDD", X"0182", X"FF80", X"FF4A", X"FE61", X"FEF8", X"FF5A", X"FF38", X"FF61", X"0203", X"010E", X"0091", X"0199", X"0351", X"03DF", X"060C", X"01CB", X"023E", X"0093", X"01F0", X"072B", X"0499", X"0307", X"0751", X"0607", X"028D", X"038B", X"049A", X"0320", X"022F", X"0169", X"001A", X"0147", X"FFBE", X"016E"),
--        (X"FF13", X"0121", X"FF94", X"FFF8", X"0049", X"0057", X"FE6D", X"0012", X"FEF7", X"FF27", X"0074", X"FF3D", X"FF38", X"FF24", X"0062", X"FFB7", X"FF0B", X"0094", X"0074", X"FF4A", X"0105", X"0029", X"FFBA", X"FFB6", X"FF90", X"FFAC", X"FFBC", X"FFDD", X"011F", X"0078", X"006C", X"FFE1", X"FFBE", X"005C", X"FCEE", X"FE01", X"FCB7", X"FDAC", X"FC5A", X"FDC9", X"FFB5", X"FE13", X"FCF0", X"FCB8", X"FF5F", X"FF02", X"FE5B", X"FBFB", X"FD53", X"FF29", X"FE1D", X"FF0F", X"FD62", X"01D4", X"007C", X"004A", X"FEA0", X"FF91", X"FFF1", X"022C", X"0034", X"00E5", X"FD55", X"FD8F", X"FC2F", X"FA98", X"F89F", X"F90E", X"F9CF", X"F9EC", X"F709", X"F849", X"F960", X"FA13", X"F95F", X"FC2D", X"FC1F", X"FB93", X"FE8B", X"FB34", X"FD7F", X"0002", X"FEA7", X"FF16", X"0080", X"FF58", X"01B9", X"0168", X"0235", X"FCE8", X"FB28", X"FB3D", X"FB9A", X"FBEC", X"FC75", X"FBB6", X"FAEF", X"FB18", X"FCD8", X"FD2F", X"FDF8", X"FDD4", X"FCA0", X"FD91", X"0029", X"FD92", X"FBAE", X"FC1C", X"FF7E", X"007D", X"00B0", X"FF13", X"FFF4", X"FF86", X"FEBD", X"00C2", X"FC81", X"F9D3", X"F884", X"FA91", X"F94F", X"FC11", X"FCFC", X"FEC5", X"FC25", X"FC1F", X"FBCC", X"FD9E", X"FE6A", X"FD36", X"FE58", X"FED8", X"FEA7", X"006C", X"00EA", X"036F", X"0322", X"015D", X"0176", X"FEB9", X"FF93", X"FFBB", X"FDDF", X"FFAF", X"F9A0", X"FAFE", X"FB41", X"FBD1", X"FE79", X"FFB0", X"0133", X"026F", X"016E", X"02BB", X"02B2", X"006A", X"FEAC", X"0066", X"0121", X"0177", X"01EF", X"0357", X"02B8", X"0326", X"01FC", X"0332", X"030D", X"FE26", X"FFEC", X"FF80", X"01B2", X"FE59", X"FEF2", X"FE77", X"FE4C", X"FF1D", X"0153", X"01A8", X"0268", X"02B6", X"0259", X"02A3", X"0388", X"00BE", X"00A1", X"0151", X"024D", X"03DF", X"0176", X"0199", X"022E", X"0162", X"00F4", X"0509", X"01F7", X"FFB4", X"FFBC", X"FDD3", X"007F", X"FF9D", X"FB30", X"FF4D", X"FE90", X"0000", X"01B4", X"0254", X"02A2", X"0227", X"0359", X"04B0", X"03B1", X"024F", X"0384", X"02E0", X"0335", X"0175", X"0377", X"0253", X"00C8", X"0021", X"FF75", X"02B8", X"00CE", X"0327", X"03D3", X"FF69", X"0284", X"FF0F", X"FB9A", X"FEF3", X"FEF6", X"0130", X"0286", X"022B", X"0181", X"033A", X"0262", X"009A", X"016A", X"0133", X"023A", X"0008", X"0237", X"FFC1", X"0239", X"008D", X"FD2F", X"FF31", X"00BD", X"FFDA", X"FF38", X"FF99", X"0049", X"01A4", X"0071", X"FFD6", X"FC5F", X"FE6B", X"001D", X"0031", X"01BD", X"FF93", X"029C", X"042B", X"032F", X"0342", X"003E", X"0182", X"0011", X"FFCE", X"00BB", X"FEAB", X"FE29", X"FDC7", X"FC2C", X"FB64", X"FEB2", X"FE4A", X"FF1E", X"0240", X"00AE", X"FEFB", X"01A7", X"003B", X"FDFF", X"015A", X"FE96", X"005E", X"0390", X"04C3", X"0450", X"058C", X"03A9", X"00C1", X"FD71", X"FE63", X"00ED", X"FE97", X"FE32", X"FDDB", X"FE98", X"FD32", X"FCE1", X"FA6C", X"FCCB", X"00A5", X"0145", X"00B3", X"FFF3", X"0282", X"0130", X"FD7B", X"FE26", X"0127", X"0345", X"038C", X"0326", X"0254", X"0483", X"05C3", X"00C0", X"FBC0", X"F8C6", X"FDBC", X"001E", X"0217", X"0168", X"FE01", X"FFC5", X"002C", X"FFB6", X"FBF1", X"FB1D", X"FCB3", X"FF31", X"FE1D", X"FFD5", X"025B", X"01FD", X"0056", X"02E0", X"0362", X"04C3", X"055D", X"02F0", X"00C5", X"0226", X"FFC7", X"FA95", X"F82D", X"F8CE", X"FB9B", X"FE55", X"00F4", X"0338", X"01D7", X"FFA9", X"FF3B", X"0154", X"00B2", X"FD10", X"FE20", X"FF0C", X"FEAB", X"FFEB", X"01E1", X"0138", X"0303", X"0612", X"03D2", X"03D1", X"051E", X"017E", X"02C9", X"0093", X"FD82", X"FC2F", X"F985", X"F853", X"FB1A", X"FC83", X"FFEB", X"0037", X"013A", X"015E", X"FFFD", X"015A", X"00BB", X"000A", X"FD09", X"FBEE", X"FD34", X"020A", X"FEAB", X"FFEB", X"034A", X"0559", X"04D8", X"03E2", X"0488", X"0189", X"0152", X"FFAE", X"FD83", X"FA19", X"F95D", X"F8A4", X"F97F", X"FCBA", X"FF57", X"00E0", X"003B", X"0290", X"020A", X"02E0", X"0400", X"031D", X"FD2F", X"FE66", X"FDF7", X"02CF", X"FE6B", X"FDDE", X"FD13", X"0379", X"0467", X"0177", X"01AA", X"0006", X"FE41", X"006B", X"FF22", X"FC65", X"F7AE", X"F57A", X"F989", X"FCA6", X"0206", X"03AF", X"013A", X"0183", X"0247", X"01CC", X"0107", X"0135", X"FCCA", X"FE19", X"FE79", X"00A3", X"FE14", X"FDEF", X"FB36", X"00B8", X"034F", X"FFA1", X"0074", X"0034", X"FFD9", X"FFCB", X"FE8C", X"FC4C", X"F65C", X"F47C", X"FB47", X"00A6", X"0283", X"0224", X"029F", X"00D4", X"FFFE", X"013A", X"003E", X"FF71", X"FC77", X"F99C", X"FDE0", X"00C4", X"FDB9", X"FBEC", X"FC4E", X"00E5", X"FFDA", X"FF8B", X"FE76", X"FED2", X"FF1F", X"01C2", X"FF4B", X"F9E9", X"F59A", X"F731", X"0165", X"043F", X"05CA", X"02F1", X"0184", X"00F3", X"015B", X"006E", X"FD06", X"FCA7", X"FDA1", X"FC52", X"0219", X"0229", X"FE69", X"FFA1", X"FC9B", X"00AB", X"FF0D", X"FDC8", X"FEA1", X"FF27", X"FE4C", X"0014", X"FE50", X"F742", X"F743", X"FE67", X"0337", X"027B", X"020B", X"00C5", X"00D3", X"009D", X"FF6C", X"FE0C", X"FC1D", X"FC93", X"FF7A", X"FE25", X"FE86", X"FFA5", X"FEF0", X"0272", X"FF98", X"01FD", X"FCC2", X"FCE6", X"FD9D", X"FDB3", X"FC92", X"FBFA", X"FD22", X"F9E0", X"FB9A", X"02A4", X"0374", X"0159", X"FF0F", X"FE89", X"FE8B", X"FDD6", X"FCA7", X"FA57", X"FB7A", X"01A7", X"FFEF", X"FD14", X"00C4", X"FFBE", X"01CC", X"01FC", X"0102", X"0176", X"0097", X"FDA6", X"FC4A", X"FCA5", X"FA34", X"FB1C", X"FBD8", X"FD0F", X"014F", X"01BB", X"0102", X"FFB1", X"FFC8", X"FEF7", X"FF1A", X"F9AA", X"FBF6", X"FAB1", X"FBD9", X"01BC", X"037C", X"FDA1", X"0002", X"0186", X"FE6B", X"FE12", X"FD5C", X"FD61", X"FE2D", X"FEC9", X"FE48", X"FBC5", X"FC97", X"FEBE", X"FF43", X"00C5", X"0171", X"0153", X"01F4", X"01C5", X"FEA1", X"FE57", X"FCDF", X"FBDA", X"FD43", X"FF11", X"FE80", X"02F7", X"052A", X"020F", X"0028", X"00E6", X"FF78", X"FEB7", X"FA0A", X"FB8C", X"FDE5", X"FD33", X"FD35", X"FE5E", X"0047", X"01BA", X"02DB", X"01B6", X"0306", X"02DE", X"020F", X"0267", X"FF87", X"FFC7", X"FD46", X"FDFE", X"FEF8", X"FE7D", X"00B4", X"05F1", X"042F", X"0244", X"FEBD", X"002C", X"FF3B", X"FAB9", X"FDDC", X"FB31", X"FE5D", X"FD6C", X"FC1D", X"FDE3", X"FE78", X"FFE8", X"0052", X"0293", X"0056", X"02BF", X"0142", X"0176", X"01A5", X"FE0B", X"FF0B", X"FD9C", X"0180", X"01A2", X"0325", X"070E", X"03BB", X"0109", X"0098", X"FEC0", X"FFF2", X"001E", X"FF0D", X"FDF9", X"0039", X"FD8D", X"FC04", X"FC14", X"FE0C", X"FE1F", X"FB25", X"FE08", X"005D", X"FF06", X"0031", X"0083", X"03BD", X"009D", X"020B", X"029D", X"0173", X"03C9", X"05ED", X"0374", X"FED5", X"FE80", X"0002", X"007B", X"00D2", X"FF4F", X"043A", X"028E", X"0031", X"0054", X"FEDC", X"FBFB", X"FC20", X"FC11", X"FD44", X"FE0C", X"FE57", X"FE99", X"FF87", X"00C9", X"0065", X"0351", X"0313", X"0284", X"0600", X"04D3", X"0334", X"0517", X"00A1", X"FF34", X"00DA", X"FE57", X"FE83", X"FFF0", X"FFF9", X"0150", X"0231", X"02BA", X"02F8", X"03E9", X"05DF", X"03EB", X"0488", X"0570", X"04E5", X"06A0", X"06E6", X"028D", X"0432", X"0395", X"04B9", X"06C6", X"069D", X"05BF", X"0271", X"0115", X"00FE", X"FF36", X"FFAF", X"00CF", X"FFA9", X"011B", X"005D", X"00DD", X"008D", X"028F", X"0415", X"0247", X"04AA", X"05ED", X"04E3", X"0584", X"0321", X"0682", X"032E", X"036C", X"0299", X"02C4", X"04A0", X"0446", X"0369", X"03CF", X"FF16", X"FFDF", X"0160", X"FFB4", X"00AD"),
--        (X"FE56", X"FF38", X"00E6", X"FFA3", X"00CC", X"FFF8", X"FFE3", X"FF93", X"00BE", X"FFCF", X"0055", X"00F8", X"FFD4", X"FFA8", X"FFFE", X"01C2", X"FFFD", X"0040", X"0124", X"FF3F", X"0097", X"FF9F", X"003E", X"FE97", X"FF27", X"00A2", X"FF5D", X"FFF0", X"015F", X"FF18", X"FF99", X"FF5A", X"0082", X"0020", X"FF2C", X"FF0E", X"00C5", X"003A", X"FDAD", X"0203", X"016F", X"0233", X"0002", X"0496", X"036D", X"01D8", X"FE3A", X"0033", X"FE14", X"FE38", X"FF23", X"FE49", X"0051", X"00C9", X"0094", X"FF6C", X"FFD7", X"00C1", X"002B", X"0335", X"02E7", X"FF0D", X"FE08", X"FD4D", X"FB4E", X"F94D", X"F886", X"FC8A", X"FE37", X"FEB3", X"FC89", X"FFF0", X"028C", X"007C", X"01D3", X"FDF0", X"FD85", X"FD80", X"FF7B", X"FE8E", X"FB8A", X"FDAE", X"0155", X"0066", X"FF91", X"0025", X"01D4", X"0297", X"FDAD", X"FC8F", X"FE9F", X"FDB6", X"02D9", X"FCCC", X"FEF0", X"0033", X"01CF", X"004E", X"0368", X"0431", X"02AD", X"039D", X"02D0", X"FF94", X"FF1F", X"FF60", X"FCCF", X"FCC3", X"FC6F", X"FF81", X"FC47", X"0000", X"0021", X"FEA6", X"039F", X"048A", X"FF3F", X"FD98", X"FD0F", X"FCB2", X"FD39", X"FC4C", X"FB09", X"FB85", X"FE44", X"01E8", X"0045", X"01A1", X"FF9B", X"FFF9", X"0051", X"FDF1", X"FDA1", X"FE3F", X"FDFF", X"FE3A", X"FECE", X"FF8C", X"02EE", X"0065", X"FFB6", X"FFF2", X"FF6E", X"FFEC", X"FBC5", X"FF22", X"FE1A", X"FD20", X"FCD3", X"FD42", X"FE11", X"FF82", X"00BF", X"019C", X"0172", X"FF6F", X"FFE4", X"FE36", X"FDD1", X"FF2D", X"006F", X"FF37", X"FF54", X"FD69", X"FDD4", X"00E6", X"0018", X"FE8C", X"FF82", X"0045", X"00C8", X"0277", X"FD83", X"000A", X"0096", X"FEF2", X"01B2", X"01FF", X"03CF", X"03E1", X"0607", X"0473", X"03B4", X"021F", X"020D", X"0251", X"0305", X"FFE2", X"024A", X"0210", X"FFFA", X"002A", X"0019", X"FFA1", X"FE92", X"FE63", X"FF8C", X"0198", X"FFA1", X"04A8", X"FE3D", X"00F4", X"FFE0", X"01FC", X"053C", X"056C", X"0729", X"03BC", X"040F", X"0411", X"035E", X"02CD", X"0344", X"057F", X"0375", X"0268", X"02FE", X"0263", X"FFDA", X"013D", X"00E6", X"011A", X"FEAC", X"FDFE", X"01F1", X"0112", X"FF17", X"0316", X"FEE3", X"00EA", X"0195", X"0478", X"06B8", X"0487", X"04BE", X"0379", X"00C5", X"028A", X"0059", X"027B", X"0438", X"0422", X"0643", X"03DB", X"0260", X"00E5", X"0260", X"0305", X"02F9", X"02A6", X"0030", X"02B0", X"FFEC", X"03F1", X"FEEF", X"01AE", X"00D7", X"0093", X"027A", X"057B", X"03F9", X"0241", X"007A", X"00CB", X"0057", X"0141", X"003D", X"01A7", X"02BD", X"0679", X"03B9", X"030F", X"02F2", X"01FF", X"024C", X"049C", X"072A", X"07AE", X"03C6", X"03DD", X"0085", X"0239", X"02EC", X"026B", X"FF5A", X"020B", X"0297", X"00DC", X"025D", X"FFA3", X"01A3", X"018A", X"018D", X"03E4", X"06A4", X"0622", X"0743", X"052F", X"0458", X"0359", X"0514", X"0186", X"0372", X"061B", X"097A", X"0874", X"07AE", X"0372", X"00B5", X"0215", X"0600", X"0167", X"00C5", X"0029", X"016F", X"003D", X"FFED", X"FE3B", X"0006", X"028E", X"040A", X"0B35", X"0B5C", X"0AA8", X"071B", X"03F6", X"02A5", X"0088", X"0244", X"011A", X"0438", X"055C", X"0810", X"089C", X"07A6", X"0328", X"0020", X"01B0", X"0474", X"0273", X"0070", X"010D", X"00F5", X"0141", X"FD6C", X"FD13", X"FEC5", X"FF8A", X"034B", X"06CE", X"07AE", X"0610", X"018D", X"011E", X"FF2D", X"FBA2", X"FF8C", X"FE46", X"0164", X"0414", X"0379", X"01C5", X"0491", X"0382", X"FF4A", X"01FA", X"0436", X"01A1", X"0110", X"FDD2", X"0009", X"FDDE", X"FE37", X"FD31", X"FB84", X"FD01", X"FF1C", X"0288", X"015F", X"FEFF", X"FDA1", X"FDE9", X"FCF8", X"FCF1", X"FE0F", X"0070", X"014F", X"013D", X"0103", X"FEA7", X"FEEF", X"FCBC", X"0141", X"0293", X"03AC", X"FE9C", X"FE89", X"FF38", X"FE84", X"F9AC", X"FCE1", X"FD49", X"FDFD", X"FA7C", X"FCE2", X"FC3C", X"FD60", X"FC4B", X"FC3D", X"FDA8", X"FFB5", X"0104", X"00EB", X"028B", X"032B", X"00B0", X"02CA", X"FF8F", X"FB25", X"FEB6", X"0045", X"028F", X"00F7", X"FEF7", X"FFC5", X"008C", X"FE4F", X"FD81", X"FCC5", X"FE22", X"FDBC", X"FCA9", X"FD63", X"FCCE", X"FB25", X"FA88", X"F9E2", X"FA59", X"FF19", X"0036", X"031B", X"02AA", X"016F", X"0347", X"02CD", X"FB1F", X"F7B5", X"FC95", X"FED6", X"027D", X"00E4", X"FF22", X"0027", X"0084", X"FD42", X"FD9D", X"FE1C", X"FF76", X"FDE7", X"FB63", X"FB4E", X"FA39", X"FBF0", X"FAF4", X"F884", X"FBC9", X"FEE7", X"FF15", X"00C9", X"FDDE", X"0009", X"0107", X"FE3C", X"F681", X"F835", X"FD5F", X"FF55", X"023A", X"FE95", X"01F4", X"0081", X"002E", X"0126", X"FC3D", X"FCD5", X"FE98", X"FDC9", X"FCBF", X"FC31", X"FB68", X"FA64", X"F98B", X"F8E6", X"FC78", X"FCDC", X"FE18", X"FEBE", X"FDC2", X"FE56", X"FF1A", X"000B", X"F99B", X"FD31", X"01EB", X"026A", X"FFC7", X"02E0", X"FF96", X"FDF2", X"FFE0", X"FC91", X"FB5A", X"FF20", X"000C", X"FFA2", X"FEFA", X"FCF3", X"FDFC", X"FCFA", X"FB71", X"FA6C", X"FD40", X"FDBC", X"FEB6", X"FF2E", X"FEF2", X"FEF2", X"FA95", X"FAA4", X"F962", X"FD7D", X"FB94", X"00A2", X"0385", X"03E4", X"FEB2", X"FE8E", X"FDDE", X"FFF9", X"FF38", X"00A3", X"022E", X"0003", X"009F", X"FFD6", X"FF54", X"FE80", X"FA8B", X"FAB5", X"FDA6", X"FEA5", X"FFE7", X"FDD5", X"FD09", X"FE02", X"FD93", X"FB96", X"FB4B", X"F9B1", X"FCEE", X"012D", X"0404", X"0320", X"FD4E", X"FD89", X"0025", X"FF94", X"0021", X"00A5", X"0385", X"01E2", X"0294", X"FFCC", X"FE9C", X"FCD1", X"FCBB", X"FD26", X"FD1C", X"FD33", X"FF27", X"FD88", X"FD3C", X"0009", X"FDE6", X"FC2A", X"F9C5", X"FD39", X"0229", X"011D", X"FE0B", X"01C9", X"012F", X"FE2C", X"0208", X"02D5", X"028D", X"FF98", X"01B8", X"004E", X"002F", X"FF3A", X"00F8", X"006B", X"FF88", X"012E", X"FF42", X"FDF7", X"FDA5", X"FD61", X"001C", X"FE20", X"FBDC", X"FC23", X"FD03", X"FD6B", X"00FA", X"002D", X"FED3", X"0013", X"FE31", X"FDC6", X"00DC", X"03FE", X"0327", X"02B2", X"0055", X"FF7F", X"00E0", X"0037", X"02D5", X"042C", X"0483", X"0228", X"0200", X"0035", X"FD3B", X"FD40", X"FC0E", X"FDB9", X"FDBE", X"FBAE", X"FDAA", X"FE80", X"010B", X"006F", X"FF52", X"FF69", X"010D", X"FF9E", X"035E", X"04E8", X"044D", X"025B", X"0285", X"0302", X"02E4", X"0424", X"0597", X"0526", X"05D8", X"060C", X"04FB", X"FF1E", X"FC3E", X"FC32", X"FC87", X"FE2D", X"FF17", X"FE6A", X"FCB7", X"FDCD", X"FF43", X"004B", X"FFAC", X"00EF", X"04D2", X"057F", X"06BD", X"04AC", X"03B7", X"02EC", X"038C", X"0476", X"044A", X"052B", X"04B9", X"049E", X"066B", X"027F", X"021E", X"FEE6", X"FDDA", X"FC8C", X"FE57", X"FBEC", X"FEE0", X"00F7", X"FC45", X"FDBE", X"FE84", X"01B4", X"FF34", X"FE33", X"0361", X"0253", X"03BD", X"003B", X"FF6B", X"027F", X"0150", X"00FE", X"0100", X"0012", X"0026", X"00BA", X"0055", X"010A", X"039B", X"02B4", X"015B", X"FC8A", X"FE15", X"FFCF", X"0133", X"0425", X"FCB3", X"FF77", X"006B", X"0079", X"00F0", X"005F", X"FF76", X"FB8A", X"FD87", X"FEAA", X"FDE0", X"FE51", X"02CB", X"0156", X"FF81", X"FE57", X"0198", X"0228", X"01EA", X"02EC", X"0366", X"0401", X"02EC", X"00DB", X"0102", X"020F", X"003A", X"031F", X"00B2", X"FFC0", X"FFB3", X"FEFD", X"008A", X"FF8D", X"011F", X"FFA1", X"0053", X"0157", X"0161", X"02A5", X"01B6", X"03A2", X"FFDC", X"FF53", X"0465", X"010A", X"0118", X"037D", X"0440", X"0151", X"008B", X"FF5F", X"021E", X"02A1", X"037A", X"FECF", X"00EB", X"FF04", X"0025")
    );
    
    

begin
    

    
   
   uut: entity work.mat_mult(Structural)
               generic map(
                           M => M,
                           N => N
               )
               
               port map( 
                         Aprev => X,
                         W => W1,
                         Z => Z
               );



end Stimulus;
