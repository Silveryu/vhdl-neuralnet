----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 05/27/2018 02:17:04 PM
-- Design Name: 
-- Module Name: normalize - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.all;


-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity normalize is
    -- N : length of input
    -- DIV : value with which to normalize
    port ( 
        dataIn : in std_logic_vector(7 downto 0);
        dataOut : out std_logic_vector(15 downto 0)
    );
end normalize;

architecture Behavioral of normalize is 
    -- decimal part : N-1, fractional part : -B
    --  ^ ufixed(N-1 downto -B)
    -- Q3.12
begin
process (dataIn) is
	begin
		case dataIn is
			when "00000000" => dataOut <= "0000000000000000";
			when "00000001" => dataOut <= "0000000000010000";
			when "00000010" => dataOut <= "0000000000100000";
			when "00000011" => dataOut <= "0000000000110000";
			when "00000100" => dataOut <= "0000000001000000";
			when "00000101" => dataOut <= "0000000001010000";
			when "00000110" => dataOut <= "0000000001100000";
			when "00000111" => dataOut <= "0000000001110000";
			when "00001000" => dataOut <= "0000000010000001";
			when "00001001" => dataOut <= "0000000010010001";
			when "00001010" => dataOut <= "0000000010100001";
			when "00001011" => dataOut <= "0000000010110001";
			when "00001100" => dataOut <= "0000000011000001";
			when "00001101" => dataOut <= "0000000011010001";
			when "00001110" => dataOut <= "0000000011100001";
			when "00001111" => dataOut <= "0000000011110001";
			when "00010000" => dataOut <= "0000000100000001";
			when "00010001" => dataOut <= "0000000100010001";
			when "00010010" => dataOut <= "0000000100100001";
			when "00010011" => dataOut <= "0000000100110001";
			when "00010100" => dataOut <= "0000000101000001";
			when "00010101" => dataOut <= "0000000101010001";
			when "00010110" => dataOut <= "0000000101100001";
			when "00010111" => dataOut <= "0000000101110001";
			when "00011000" => dataOut <= "0000000110000010";
			when "00011001" => dataOut <= "0000000110010010";
			when "00011010" => dataOut <= "0000000110100010";
			when "00011011" => dataOut <= "0000000110110010";
			when "00011100" => dataOut <= "0000000111000010";
			when "00011101" => dataOut <= "0000000111010010";
			when "00011110" => dataOut <= "0000000111100010";
			when "00011111" => dataOut <= "0000000111110010";
			when "00100000" => dataOut <= "0000001000000010";
			when "00100001" => dataOut <= "0000001000010010";
			when "00100010" => dataOut <= "0000001000100010";
			when "00100011" => dataOut <= "0000001000110010";
			when "00100100" => dataOut <= "0000001001000010";
			when "00100101" => dataOut <= "0000001001010010";
			when "00100110" => dataOut <= "0000001001100010";
			when "00100111" => dataOut <= "0000001001110010";
			when "00101000" => dataOut <= "0000001010000011";
			when "00101001" => dataOut <= "0000001010010011";
			when "00101010" => dataOut <= "0000001010100011";
			when "00101011" => dataOut <= "0000001010110011";
			when "00101100" => dataOut <= "0000001011000011";
			when "00101101" => dataOut <= "0000001011010011";
			when "00101110" => dataOut <= "0000001011100011";
			when "00101111" => dataOut <= "0000001011110011";
			when "00110000" => dataOut <= "0000001100000011";
			when "00110001" => dataOut <= "0000001100010011";
			when "00110010" => dataOut <= "0000001100100011";
			when "00110011" => dataOut <= "0000001100110011";
			when "00110100" => dataOut <= "0000001101000011";
			when "00110101" => dataOut <= "0000001101010011";
			when "00110110" => dataOut <= "0000001101100011";
			when "00110111" => dataOut <= "0000001101110011";
			when "00111000" => dataOut <= "0000001110000100";
			when "00111001" => dataOut <= "0000001110010100";
			when "00111010" => dataOut <= "0000001110100100";
			when "00111011" => dataOut <= "0000001110110100";
			when "00111100" => dataOut <= "0000001111000100";
			when "00111101" => dataOut <= "0000001111010100";
			when "00111110" => dataOut <= "0000001111100100";
			when "00111111" => dataOut <= "0000001111110100";
			when "01000000" => dataOut <= "0000010000000100";
			when "01000001" => dataOut <= "0000010000010100";
			when "01000010" => dataOut <= "0000010000100100";
			when "01000011" => dataOut <= "0000010000110100";
			when "01000100" => dataOut <= "0000010001000100";
			when "01000101" => dataOut <= "0000010001010100";
			when "01000110" => dataOut <= "0000010001100100";
			when "01000111" => dataOut <= "0000010001110100";
			when "01001000" => dataOut <= "0000010010000101";
			when "01001001" => dataOut <= "0000010010010101";
			when "01001010" => dataOut <= "0000010010100101";
			when "01001011" => dataOut <= "0000010010110101";
			when "01001100" => dataOut <= "0000010011000101";
			when "01001101" => dataOut <= "0000010011010101";
			when "01001110" => dataOut <= "0000010011100101";
			when "01001111" => dataOut <= "0000010011110101";
			when "01010000" => dataOut <= "0000010100000101";
			when "01010001" => dataOut <= "0000010100010101";
			when "01010010" => dataOut <= "0000010100100101";
			when "01010011" => dataOut <= "0000010100110101";
			when "01010100" => dataOut <= "0000010101000101";
			when "01010101" => dataOut <= "0000010101010101";
			when "01010110" => dataOut <= "0000010101100101";
			when "01010111" => dataOut <= "0000010101110101";
			when "01011000" => dataOut <= "0000010110000110";
			when "01011001" => dataOut <= "0000010110010110";
			when "01011010" => dataOut <= "0000010110100110";
			when "01011011" => dataOut <= "0000010110110110";
			when "01011100" => dataOut <= "0000010111000110";
			when "01011101" => dataOut <= "0000010111010110";
			when "01011110" => dataOut <= "0000010111100110";
			when "01011111" => dataOut <= "0000010111110110";
			when "01100000" => dataOut <= "0000011000000110";
			when "01100001" => dataOut <= "0000011000010110";
			when "01100010" => dataOut <= "0000011000100110";
			when "01100011" => dataOut <= "0000011000110110";
			when "01100100" => dataOut <= "0000011001000110";
			when "01100101" => dataOut <= "0000011001010110";
			when "01100110" => dataOut <= "0000011001100110";
			when "01100111" => dataOut <= "0000011001110110";
			when "01101000" => dataOut <= "0000011010000111";
			when "01101001" => dataOut <= "0000011010010111";
			when "01101010" => dataOut <= "0000011010100111";
			when "01101011" => dataOut <= "0000011010110111";
			when "01101100" => dataOut <= "0000011011000111";
			when "01101101" => dataOut <= "0000011011010111";
			when "01101110" => dataOut <= "0000011011100111";
			when "01101111" => dataOut <= "0000011011110111";
			when "01110000" => dataOut <= "0000011100000111";
			when "01110001" => dataOut <= "0000011100010111";
			when "01110010" => dataOut <= "0000011100100111";
			when "01110011" => dataOut <= "0000011100110111";
			when "01110100" => dataOut <= "0000011101000111";
			when "01110101" => dataOut <= "0000011101010111";
			when "01110110" => dataOut <= "0000011101100111";
			when "01110111" => dataOut <= "0000011101110111";
			when "01111000" => dataOut <= "0000011110001000";
			when "01111001" => dataOut <= "0000011110011000";
			when "01111010" => dataOut <= "0000011110101000";
			when "01111011" => dataOut <= "0000011110111000";
			when "01111100" => dataOut <= "0000011111001000";
			when "01111101" => dataOut <= "0000011111011000";
			when "01111110" => dataOut <= "0000011111101000";
			when "01111111" => dataOut <= "0000011111111000";
			when "10000000" => dataOut <= "0000100000001000";
			when "10000001" => dataOut <= "0000100000011000";
			when "10000010" => dataOut <= "0000100000101000";
			when "10000011" => dataOut <= "0000100000111000";
			when "10000100" => dataOut <= "0000100001001000";
			when "10000101" => dataOut <= "0000100001011000";
			when "10000110" => dataOut <= "0000100001101000";
			when "10000111" => dataOut <= "0000100001111000";
			when "10001000" => dataOut <= "0000100010001001";
			when "10001001" => dataOut <= "0000100010011001";
			when "10001010" => dataOut <= "0000100010101001";
			when "10001011" => dataOut <= "0000100010111001";
			when "10001100" => dataOut <= "0000100011001001";
			when "10001101" => dataOut <= "0000100011011001";
			when "10001110" => dataOut <= "0000100011101001";
			when "10001111" => dataOut <= "0000100011111001";
			when "10010000" => dataOut <= "0000100100001001";
			when "10010001" => dataOut <= "0000100100011001";
			when "10010010" => dataOut <= "0000100100101001";
			when "10010011" => dataOut <= "0000100100111001";
			when "10010100" => dataOut <= "0000100101001001";
			when "10010101" => dataOut <= "0000100101011001";
			when "10010110" => dataOut <= "0000100101101001";
			when "10010111" => dataOut <= "0000100101111001";
			when "10011000" => dataOut <= "0000100110001010";
			when "10011001" => dataOut <= "0000100110011010";
			when "10011010" => dataOut <= "0000100110101010";
			when "10011011" => dataOut <= "0000100110111010";
			when "10011100" => dataOut <= "0000100111001010";
			when "10011101" => dataOut <= "0000100111011010";
			when "10011110" => dataOut <= "0000100111101010";
			when "10011111" => dataOut <= "0000100111111010";
			when "10100000" => dataOut <= "0000101000001010";
			when "10100001" => dataOut <= "0000101000011010";
			when "10100010" => dataOut <= "0000101000101010";
			when "10100011" => dataOut <= "0000101000111010";
			when "10100100" => dataOut <= "0000101001001010";
			when "10100101" => dataOut <= "0000101001011010";
			when "10100110" => dataOut <= "0000101001101010";
			when "10100111" => dataOut <= "0000101001111010";
			when "10101000" => dataOut <= "0000101010001011";
			when "10101001" => dataOut <= "0000101010011011";
			when "10101010" => dataOut <= "0000101010101011";
			when "10101011" => dataOut <= "0000101010111011";
			when "10101100" => dataOut <= "0000101011001011";
			when "10101101" => dataOut <= "0000101011011011";
			when "10101110" => dataOut <= "0000101011101011";
			when "10101111" => dataOut <= "0000101011111011";
			when "10110000" => dataOut <= "0000101100001011";
			when "10110001" => dataOut <= "0000101100011011";
			when "10110010" => dataOut <= "0000101100101011";
			when "10110011" => dataOut <= "0000101100111011";
			when "10110100" => dataOut <= "0000101101001011";
			when "10110101" => dataOut <= "0000101101011011";
			when "10110110" => dataOut <= "0000101101101011";
			when "10110111" => dataOut <= "0000101101111011";
			when "10111000" => dataOut <= "0000101110001100";
			when "10111001" => dataOut <= "0000101110011100";
			when "10111010" => dataOut <= "0000101110101100";
			when "10111011" => dataOut <= "0000101110111100";
			when "10111100" => dataOut <= "0000101111001100";
			when "10111101" => dataOut <= "0000101111011100";
			when "10111110" => dataOut <= "0000101111101100";
			when "10111111" => dataOut <= "0000101111111100";
			when "11000000" => dataOut <= "0000110000001100";
			when "11000001" => dataOut <= "0000110000011100";
			when "11000010" => dataOut <= "0000110000101100";
			when "11000011" => dataOut <= "0000110000111100";
			when "11000100" => dataOut <= "0000110001001100";
			when "11000101" => dataOut <= "0000110001011100";
			when "11000110" => dataOut <= "0000110001101100";
			when "11000111" => dataOut <= "0000110001111100";
			when "11001000" => dataOut <= "0000110010001101";
			when "11001001" => dataOut <= "0000110010011101";
			when "11001010" => dataOut <= "0000110010101101";
			when "11001011" => dataOut <= "0000110010111101";
			when "11001100" => dataOut <= "0000110011001101";
			when "11001101" => dataOut <= "0000110011011101";
			when "11001110" => dataOut <= "0000110011101101";
			when "11001111" => dataOut <= "0000110011111101";
			when "11010000" => dataOut <= "0000110100001101";
			when "11010001" => dataOut <= "0000110100011101";
			when "11010010" => dataOut <= "0000110100101101";
			when "11010011" => dataOut <= "0000110100111101";
			when "11010100" => dataOut <= "0000110101001101";
			when "11010101" => dataOut <= "0000110101011101";
			when "11010110" => dataOut <= "0000110101101101";
			when "11010111" => dataOut <= "0000110101111101";
			when "11011000" => dataOut <= "0000110110001110";
			when "11011001" => dataOut <= "0000110110011110";
			when "11011010" => dataOut <= "0000110110101110";
			when "11011011" => dataOut <= "0000110110111110";
			when "11011100" => dataOut <= "0000110111001110";
			when "11011101" => dataOut <= "0000110111011110";
			when "11011110" => dataOut <= "0000110111101110";
			when "11011111" => dataOut <= "0000110111111110";
			when "11100000" => dataOut <= "0000111000001110";
			when "11100001" => dataOut <= "0000111000011110";
			when "11100010" => dataOut <= "0000111000101110";
			when "11100011" => dataOut <= "0000111000111110";
			when "11100100" => dataOut <= "0000111001001110";
			when "11100101" => dataOut <= "0000111001011110";
			when "11100110" => dataOut <= "0000111001101110";
			when "11100111" => dataOut <= "0000111001111110";
			when "11101000" => dataOut <= "0000111010001111";
			when "11101001" => dataOut <= "0000111010011111";
			when "11101010" => dataOut <= "0000111010101111";
			when "11101011" => dataOut <= "0000111010111111";
			when "11101100" => dataOut <= "0000111011001111";
			when "11101101" => dataOut <= "0000111011011111";
			when "11101110" => dataOut <= "0000111011101111";
			when "11101111" => dataOut <= "0000111011111111";
			when "11110000" => dataOut <= "0000111100001111";
			when "11110001" => dataOut <= "0000111100011111";
			when "11110010" => dataOut <= "0000111100101111";
			when "11110011" => dataOut <= "0000111100111111";
			when "11110100" => dataOut <= "0000111101001111";
			when "11110101" => dataOut <= "0000111101011111";
			when "11110110" => dataOut <= "0000111101101111";
			when "11110111" => dataOut <= "0000111101111111";
			when "11111000" => dataOut <= "0000111110010000";
			when "11111001" => dataOut <= "0000111110100000";
			when "11111010" => dataOut <= "0000111110110000";
			when "11111011" => dataOut <= "0000111111000000";
			when "11111100" => dataOut <= "0000111111010000";
			when "11111101" => dataOut <= "0000111111100000";
			when "11111110" => dataOut <= "0000111111110000";
			when others => dataOut <= "0001000000000000";
	end case;
end process;
    

end Behavioral;
