----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 05/31/2018 02:49:06 PM
-- Design Name: 
-- Module Name: weight_unit_tb - Stimulus
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;


library work;
use work.custom_type.all;


entity feed_forward_unit_tb is
end feed_forward_unit_tb;

architecture Stimulus of feed_forward_unit_tb is

    

    constant TIME_DELTA: time := 10 ns; -- clock wait time in ns
    
    constant unit_num1  : positive := 50;
    constant input_dim1 : positive := 784;
    
     constant unit_num2  : positive := 10;
     constant input_dim2 : positive := 50;

    signal X : WORD_ARRAY(0 to input_dim1-1) := (X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0030", X"0121", X"0121", X"0121", X"07E8", X"0889", X"0AFB", X"01A2", X"0A6A", X"1000", X"0F7F", X"07F8", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"01E2", X"0242", X"05E6", X"09AA", X"0AAB", X"0FE0", X"0FE0", X"0FE0", X"0FE0", X"0FE0", X"0E1E", X"0ACB", X"0FE0", X"0F2F", X"0C3C", X"0404", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0313", X"0EEF", X"0FE0", X"0FE0", X"0FE0", X"0FE0", X"0FE0", X"0FE0", X"0FE0", X"0FE0", X"0FC0", X"05D6", X"0525", X"0525", X"0384", X"0272", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0121", X"0DBE", X"0FE0", X"0FE0", X"0FE0", X"0FE0", X"0FE0", X"0C6C", X"0B6B", X"0F7F", X"0F1F", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0505", X"09CA", X"06B7", X"0FE0", X"0FE0", X"0CDD", X"00B1", X"0000", X"02B3", X"09AA", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"00E1", X"0010", X"09AA", X"0FE0", X"05A6", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"08B9", X"0FE0", X"0BEC", X"0020", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"00B1", X"0BEC", X"0FE0", X"0464", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0232", X"0F1F", X"0E1E", X"0A0A", X"06C7", X"0010", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0515", X"0F0F", X"0FE0", X"0FE0", X"0777", X"0192", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"02D3", X"0BAC", X"0FE0", X"0FE0", X"0969", X"01B2", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0101", X"05D6", X"0FD0", X"0FE0", X"0BBC", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0FA0", X"0FE0", X"0FA0", X"0404", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"02E3", X"0828", X"0B7B", X"0FE0", X"0FE0", X"0CFD", X"0020", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0272", X"0949", X"0E5E", X"0FE0", X"0FE0", X"0FE0", X"0FB0", X"0B6B", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0182", X"0727", X"0DDE", X"0FE0", X"0FE0", X"0FE0", X"0FE0", X"0C9D", X"04E5", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0171", X"0424", X"0D5D", X"0FE0", X"0FE0", X"0FE0", X"0FE0", X"0C6C", X"0515", X"0020", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0121", X"0ABB", X"0DBE", X"0FE0", X"0FE0", X"0FE0", X"0FE0", X"0C3C", X"0505", X"0091", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0373", X"0ACB", X"0E2E", X"0FE0", X"0FE0", X"0FE0", X"0FE0", X"0F4F", X"0858", X"00B1", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0889", X"0FE0", X"0FE0", X"0FE0", X"0D4D", X"0878", X"0848", X"0101", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000");    
    
    signal W1 : WORD_MAT(0 to unit_num1-1, 0 to input_dim1-1) := (	
        (X"011A", X"FF11", X"FED9", X"FFBC", X"0113", X"FF8D", X"FF6F", X"00FB", X"004E", X"004A", X"01E0", X"FF64", X"0185", X"01CB", X"FE72", X"FF2D", X"006A", X"004B", X"0088", X"0123", X"FF65", X"0135", X"FFB0", X"00DA", X"0036", X"0148", X"00F3", X"00C6", X"000A", X"FEBB", X"00D3", X"0172", X"00B8", X"00A5", X"0263", X"03C2", X"036D", X"028C", X"0534", X"0450", X"0519", X"02F0", X"00B9", X"0002", X"FC81", X"FE2C", X"0420", X"0388", X"04F4", X"04D7", X"0306", X"FFA6", X"FFF2", X"FFF7", X"FFA0", X"FF57", X"012F", X"00D5", X"000B", X"FFE9", X"02EC", X"02CE", X"0586", X"050B", X"02CE", X"0237", X"078C", X"063F", X"04EE", X"036F", X"032B", X"031F", X"0466", X"0417", X"0708", X"081C", X"04C0", X"0487", X"057F", X"053E", X"0082", X"FF38", X"FF77", X"FFFF", X"017B", X"FECB", X"FF8D", X"0080", X"0160", X"FCF0", X"FD9D", X"FAC2", X"FA87", X"F8F8", X"FA8B", X"FA62", X"FB63", X"FF5C", X"FF01", X"FEAC", X"FD3D", X"FEFB", X"01D2", X"FFD3", X"FFF4", X"00C9", X"053F", X"022C", X"FCC3", X"FBD5", X"0197", X"FF89", X"FF04", X"FD7C", X"FDDD", X"FD54", X"F9EF", X"F94D", X"FAD6", X"FAF4", X"F74A", X"FA44", X"FD9F", X"FBF1", X"FDAE", X"FC0B", X"FEF4", X"FFCD", X"FFAC", X"FF0A", X"FEFD", X"FEA3", X"016B", X"020B", X"025D", X"03D3", X"FFB4", X"FEEB", X"0257", X"FFB1", X"013C", X"FFB8", X"01D3", X"FB96", X"F598", X"F5B3", X"F682", X"F7CA", X"F991", X"F966", X"FC0C", X"FEDE", X"00A7", X"FC6E", X"FE4B", X"FDE2", X"FC50", X"FD84", X"FCF6", X"FF58", X"0162", X"FFAB", X"018E", X"0494", X"02A6", X"04D3", X"061E", X"0122", X"00E1", X"FF29", X"FE46", X"F8B9", X"F535", X"F575", X"F568", X"F83D", X"FB73", X"FCAD", X"FD46", X"FE5C", X"FF63", X"FDB5", X"FFA7", X"FF0C", X"FEBD", X"FD9A", X"FD86", X"00FA", X"FFA9", X"FF0E", X"FF61", X"03D8", X"081C", X"09DA", X"0742", X"0447", X"FDEC", X"FCA7", X"FC8D", X"F5CF", X"F3FD", X"F2EF", X"F747", X"FACA", X"FF13", X"FDC1", X"FDF9", X"FEAD", X"FEC6", X"FE30", X"0020", X"FFC8", X"FF81", X"FD48", X"FEA8", X"FE2D", X"00A0", X"01D1", X"01CF", X"0293", X"08CE", X"0AAE", X"081D", X"02C4", X"FD97", X"FC9C", X"FA43", X"F745", X"F1C8", X"F4AD", X"F8B4", X"FC85", X"FF1D", X"00AD", X"FE0D", X"FF9E", X"FF27", X"FEEB", X"FC62", X"FD45", X"FB1B", X"FC39", X"FD27", X"FD67", X"FE9A", X"0102", X"FF7A", X"032C", X"0AA4", X"0C7A", X"089F", X"0303", X"FEB6", X"FE4E", X"FAA5", X"F63A", X"F34A", X"F4D0", X"FB59", X"FF60", X"0427", X"026C", X"03F5", X"05E1", X"03AE", X"FEA0", X"FB68", X"F8EC", X"F76E", X"F878", X"F9BF", X"FBD3", X"FD83", X"00C7", X"00ED", X"038A", X"09A1", X"0A65", X"0A93", X"0389", X"FEB5", X"FEC0", X"F6EB", X"F40E", X"F4C6", X"F66B", X"FF4D", X"0763", X"08CC", X"0A31", X"0937", X"0725", X"06BA", X"02C3", X"0070", X"FCE6", X"F725", X"F64C", X"F933", X"F967", X"FB0F", X"FBFF", X"FD6A", X"0332", X"0806", X"0B06", X"0952", X"016B", X"FEA6", X"FB11", X"F895", X"F2BC", X"F3D4", X"FCFB", X"05EB", X"0B8E", X"0C2C", X"0951", X"066B", X"04D2", X"056F", X"083D", X"0960", X"05BF", X"FDB5", X"F906", X"FA11", X"FB79", X"F92E", X"FA37", X"FBD8", X"FF29", X"03D0", X"08A1", X"090E", X"017A", X"FF60", X"FBF1", X"F98E", X"F4E3", X"F6CF", X"FF0B", X"0782", X"099F", X"069B", X"0343", X"0252", X"02EF", X"0383", X"0A46", X"0BBC", X"0811", X"FFCD", X"FD14", X"FF1C", X"00D7", X"01E9", X"0044", X"FA1E", X"FABF", X"FA63", X"FF47", X"0259", X"FFBF", X"FFF6", X"FDBA", X"FA40", X"F5FF", X"F6B3", X"FDB7", X"007A", X"05FC", X"02AD", X"026F", X"021E", X"0164", X"0382", X"078E", X"0914", X"07DE", X"02CE", X"FE8F", X"015E", X"050C", X"0504", X"02F0", X"FCFF", X"F7F0", X"F6F5", X"F8A4", X"FC97", X"FDC0", X"02EE", X"FFC3", X"FC74", X"F7DD", X"F6FE", X"FC78", X"FF51", X"FE22", X"0082", X"01DE", X"0139", X"01ED", X"0373", X"069F", X"06E9", X"05EB", X"0342", X"FDF0", X"FF5A", X"FF5A", X"01B5", X"0155", X"FE41", X"F8D4", X"F7A4", X"F6A0", X"F7D6", X"FDDD", X"01CF", X"FF3C", X"FDBF", X"F889", X"F929", X"FA0D", X"F9BF", X"FB8D", X"FD7E", X"01B3", X"01C5", X"0321", X"03F6", X"07CD", X"04E8", X"042B", X"00CE", X"FED2", X"FED4", X"FD47", X"FB0B", X"FBF3", X"FAF8", X"F8BF", X"F793", X"F736", X"F77B", X"FD4E", X"FD6F", X"FEF3", X"FDEA", X"FBB3", X"FBF9", X"FBF0", X"F9C8", X"FB13", X"FECD", X"0074", X"0263", X"0261", X"02D8", X"02F9", X"03D3", X"0013", X"FE8E", X"FB6E", X"FAE0", X"FA3F", X"FAE3", X"FBE1", X"FC76", X"FE6C", X"FB83", X"F898", X"F703", X"FBD8", X"FF10", X"FF38", X"FC0A", X"FBBB", X"FD7A", X"FD94", X"FD24", X"FD1A", X"FD71", X"0069", X"02D7", X"045C", X"0330", X"048E", X"0221", X"FEBC", X"FD68", X"FACC", X"FC99", X"FBA0", X"FDC6", X"FE0A", X"FEC9", X"FF99", X"0139", X"FB1F", X"F5A3", X"FB6F", X"FF89", X"FFF1", X"F90C", X"FB0E", X"FC6A", X"FF62", X"00F6", X"FFBB", X"FF50", X"0117", X"03CA", X"04D4", X"030D", X"029F", X"0101", X"FF1D", X"FB6D", X"FB50", X"FB91", X"FC5A", X"00A1", X"FE31", X"0060", X"020A", X"042A", X"FE38", X"F863", X"FC6B", X"FECC", X"FAD0", X"FB47", X"F806", X"FAFE", X"FEB0", X"FF42", X"FE42", X"0067", X"FF2C", X"00D9", X"00BA", X"00CA", X"004C", X"FDE0", X"FE67", X"FDCF", X"FD4B", X"FD0F", X"FE15", X"0009", X"FEE2", X"00D5", X"0574", X"061C", X"FF00", X"F896", X"FC56", X"FFC0", X"FDFB", X"FB7C", X"F833", X"FA5C", X"FFB0", X"FF63", X"FF39", X"FFD5", X"FD00", X"FE28", X"FEBA", X"FED1", X"FFB0", X"FE44", X"FE83", X"FEB8", X"FF31", X"FD12", X"FD9D", X"FF56", X"FF88", X"04EC", X"0513", X"02F6", X"015C", X"FB6D", X"001A", X"00EC", X"FF50", X"FAFA", X"FB72", X"FC71", X"FFD2", X"FF37", X"FF80", X"015A", X"010B", X"FF7B", X"FE7B", X"FE9B", X"FF74", X"00CC", X"00F9", X"FECC", X"FCFE", X"FC62", X"FC6A", X"0116", X"03DF", X"02E1", X"00FF", X"00B1", X"FE8A", X"FC87", X"FD6D", X"0168", X"0050", X"FBE8", X"FB72", X"00E9", X"0129", X"FEFA", X"FEFF", X"FF64", X"FF2E", X"FF17", X"FF62", X"00AD", X"00A8", X"FF85", X"FFA7", X"00F6", X"0000", X"FE78", X"FE1F", X"FEC8", X"02CD", X"FFF0", X"0265", X"FFF1", X"FF43", X"0219", X"FF3A", X"FF4B", X"00AF", X"FE45", X"FB52", X"FDBC", X"FE7E", X"FF87", X"FDC6", X"0115", X"003C", X"FF8F", X"FE83", X"0006", X"FFF9", X"FF13", X"00A3", X"01A3", X"0130", X"FDD0", X"FCA0", X"FF84", X"FD26", X"FE73", X"01BF", X"00C0", X"FFCB", X"01BC", X"00B3", X"FF34", X"FF10", X"FF9C", X"FC71", X"F897", X"FBDA", X"FD51", X"FD51", X"FF4C", X"00D0", X"00DC", X"FEA1", X"FD1F", X"FED7", X"FC32", X"FF1C", X"0040", X"FE3F", X"015D", X"0239", X"00D3", X"FF6F", X"FE5C", X"03F7", X"00FA", X"FC11", X"FE85", X"0057", X"FF73", X"FF65", X"0229", X"013E", X"FC44", X"FA0E", X"FBAF", X"FB81", X"FACB", X"FBF8", X"FF36", X"0009", X"0009", X"0042", X"0120", X"009E", X"0356", X"046F", X"049E", X"02ED", X"03CA", X"0330", X"0480", X"083F", X"061E", X"FEF0", X"FDF1", X"FFF1", X"001F", X"FFA2", X"0013", X"00A6", X"03C6", X"FD93", X"FDE5", X"FBFF", X"FCCA", X"FDD3", X"001F", X"01AF", X"02C6", X"00D2", X"0029", X"FCC2", X"FBB6", X"FE47", X"FF8D", X"0004", X"01B3", X"FF7D", X"FD6A", X"004E", X"0224", X"FF99", X"FF47", X"FF24", X"0088", X"0016", X"FF65", X"FF13", X"004B", X"FE0A", X"00F0", X"0058", X"FEC2", X"FEAC", X"003B", X"0073", X"0059", X"F7CE", X"FD9B", X"FDE1", X"F78F", X"FB9F", X"FF01", X"FD52", X"FF6D", X"0004", X"FDD8", X"FBB5", X"FF88", X"FDB0", X"0001", X"FFF5"),
        (X"006F", X"FF68", X"00AC", X"0045", X"FFB2", X"FFF7", X"FF67", X"00BA", X"0058", X"001B", X"FF89", X"00BB", X"009A", X"00DF", X"00F4", X"007D", X"006C", X"FF1B", X"007D", X"FF4B", X"0007", X"FEB5", X"FF6F", X"009F", X"FFA8", X"0043", X"0053", X"FFC3", X"FFA3", X"0049", X"FFD0", X"FF7B", X"FEDB", X"FFB6", X"FEEC", X"00B0", X"0023", X"00EE", X"015E", X"FFA7", X"FE43", X"0209", X"FFC2", X"FF12", X"020F", X"0210", X"00D1", X"FFAD", X"0098", X"FE9D", X"FF2F", X"FE26", X"FF51", X"0071", X"010C", X"FF04", X"FF8F", X"0018", X"FF7C", X"00D1", X"00EC", X"0140", X"012A", X"00F0", X"0199", X"0482", X"05E4", X"0516", X"01E3", X"0570", X"04DD", X"0160", X"01EA", X"01B4", X"004C", X"FE7C", X"0046", X"0003", X"016B", X"0257", X"0423", X"03C5", X"FEE4", X"002E", X"FEEB", X"FF4F", X"FCAF", X"FE71", X"FF41", X"FE9D", X"0090", X"FFBD", X"0271", X"03DA", X"032C", X"02A4", X"016A", X"0276", X"01A9", X"0203", X"0133", X"00F8", X"FF31", X"FECE", X"FF73", X"FE90", X"0120", X"00E8", X"028C", X"022B", X"0040", X"FF73", X"0047", X"0005", X"FD76", X"FC58", X"FC51", X"FE45", X"FE23", X"FFF5", X"02FA", X"0555", X"04A8", X"0230", X"0292", X"00B6", X"0086", X"00A0", X"00D3", X"025E", X"00EA", X"0160", X"005B", X"FD06", X"FCF3", X"FB67", X"FDD1", X"FF62", X"FD79", X"0142", X"0021", X"FF1E", X"FEB2", X"FFB7", X"FFA4", X"FD6A", X"FDA4", X"01DF", X"04BE", X"03F5", X"0547", X"03CF", X"034A", X"012D", X"FF94", X"00EF", X"01D3", X"007D", X"FF1F", X"FD52", X"FEE4", X"004C", X"FE38", X"FD40", X"FCDC", X"FDD2", X"FC53", X"0061", X"FF0F", X"00C2", X"00F4", X"0114", X"00BE", X"0010", X"0247", X"02E5", X"048D", X"0488", X"03A4", X"01FF", X"01E2", X"000C", X"010F", X"015C", X"00D1", X"FF33", X"FF0B", X"FDD0", X"FCF6", X"FFD9", X"FFCC", X"FC1F", X"FA3D", X"FB0C", X"FCC0", X"FE67", X"0056", X"FFD2", X"049F", X"050F", X"018D", X"015D", X"032E", X"00F0", X"05FC", X"0471", X"02AD", X"01F5", X"0139", X"024C", X"FF06", X"FF29", X"FEA2", X"FEDE", X"FD37", X"FD50", X"FE2A", X"0194", X"FFC2", X"FD98", X"FB7B", X"F992", X"FC6D", X"FCEB", X"FE37", X"042D", X"0368", X"0321", X"0129", X"027B", X"01BE", X"0311", X"04AD", X"038A", X"01B9", X"014B", X"0102", X"0189", X"FED0", X"FF6F", X"FD84", X"FE50", X"FE2C", X"FE27", X"FD8F", X"FE5A", X"FE1A", X"FE38", X"F8E4", X"F8C6", X"FA8D", X"FD05", X"0217", X"0442", X"053A", X"0358", X"FF1C", X"0155", X"0274", X"02C2", X"00BC", X"0219", X"0030", X"0215", X"016F", X"FDF1", X"FE1C", X"FE09", X"FE9A", X"FF4E", X"FEAE", X"FE96", X"FE74", X"FE92", X"FC8A", X"FB97", X"F8E5", X"F848", X"F972", X"0081", X"0127", X"0255", X"0380", X"FFA7", X"0059", X"01BE", X"0323", X"0498", X"0339", X"029B", X"02D1", X"01DD", X"FE3C", X"FA56", X"F89F", X"FAE5", X"FD28", X"FEA3", X"FF3B", X"0036", X"0007", X"FFEB", X"FCD7", X"FA35", X"F53C", X"F686", X"F98B", X"0169", X"0113", X"055C", X"046D", X"0122", X"01F4", X"0466", X"03E6", X"0529", X"0449", X"05B1", X"041F", X"FDFE", X"FA9F", X"F588", X"F5FF", X"FA58", X"FBD3", X"FDDA", X"FE8F", X"013D", X"0061", X"037C", X"04A4", X"FF17", X"F82E", X"F516", X"F98B", X"FF9E", X"0116", X"048F", X"078B", X"057D", X"000B", X"04E5", X"0617", X"06C8", X"0664", X"04AC", X"01A2", X"FF12", X"F85A", X"F5D1", X"F63B", X"FBA2", X"FE31", X"FEA9", X"FFB4", X"01E5", X"0430", X"07FF", X"0C53", X"0C5F", X"0937", X"0058", X"FEA7", X"028B", X"0029", X"02BB", X"075F", X"02C3", X"FFC6", X"0448", X"06FF", X"0A14", X"0618", X"04E2", X"03F6", X"01D5", X"FA56", X"F7F5", X"FAB7", X"FBA0", X"FF80", X"0248", X"051C", X"04C9", X"0501", X"079C", X"0DD6", X"1030", X"0D7F", X"069C", X"0562", X"02EE", X"FEA2", X"FED7", X"02B9", X"00CA", X"011B", X"04C8", X"08D6", X"098E", X"0640", X"0651", X"040B", X"0047", X"F9ED", X"F9DD", X"FD47", X"01BF", X"0169", X"024D", X"04FB", X"0455", X"0369", X"03CE", X"0933", X"0BAB", X"096E", X"07AF", X"0486", X"00C0", X"FF54", X"FDAE", X"FD6C", X"006A", X"007E", X"0632", X"0745", X"0631", X"05E0", X"05A0", X"026A", X"00A8", X"FCA6", X"FF81", X"02E9", X"04C5", X"0354", X"04F1", X"0287", X"0025", X"0032", X"02E2", X"042E", X"09A6", X"0994", X"0763", X"0657", X"0270", X"0089", X"FC74", X"FD84", X"00AE", X"FC8C", X"00C1", X"0283", X"053C", X"0615", X"0517", X"043C", X"033F", X"03D7", X"0524", X"02BC", X"0201", X"0297", X"01B2", X"FEC1", X"FDA8", X"FEE6", X"FF95", X"03A7", X"083B", X"0711", X"0964", X"0451", X"031E", X"0048", X"FDF6", X"FE56", X"FB24", X"FD02", X"FF11", X"FF07", X"012E", X"017E", X"045E", X"06D6", X"0A89", X"0BAF", X"0710", X"024F", X"009D", X"FF22", X"FF9F", X"FD67", X"FDE8", X"FDED", X"FF26", X"0444", X"06AF", X"0A44", X"0863", X"055C", X"FDD6", X"01A7", X"FFFD", X"FFD3", X"FD36", X"FECA", X"FCEF", X"FA83", X"FD76", X"FED2", X"027F", X"05F5", X"07CB", X"0824", X"05F3", X"0196", X"FEF7", X"FE8E", X"FD95", X"FC3C", X"FCFE", X"FED6", X"019B", X"04EE", X"0A5A", X"09FE", X"043E", X"0308", X"FF93", X"FEE0", X"0021", X"FF5B", X"FBEB", X"FD34", X"FD30", X"FBD7", X"FC90", X"FB0A", X"FEFE", X"03D7", X"0490", X"0738", X"01DA", X"FFC9", X"FEC2", X"FF1E", X"FD25", X"FC19", X"FF13", X"00A0", X"0437", X"06D9", X"07E9", X"0569", X"0273", X"0276", X"003D", X"FF3C", X"FCA4", X"FFEA", X"FE75", X"0017", X"FE56", X"FC76", X"FBD7", X"FA45", X"FB0D", X"FE4C", X"034E", X"0407", X"02BB", X"01B5", X"00BD", X"FD32", X"FADB", X"FCFC", X"FF30", X"01FB", X"0442", X"0841", X"0952", X"046A", X"03AC", X"00B4", X"FE64", X"FDDE", X"FF20", X"FF6C", X"FF5B", X"FF20", X"FF1D", X"FC73", X"FD2D", X"FA82", X"FCB4", X"FC41", X"FF00", X"0116", X"0348", X"0237", X"FDFE", X"FE69", X"FF22", X"FECA", X"0013", X"0062", X"03A9", X"0893", X"09CF", X"0398", X"0436", X"007E", X"00AB", X"FFD2", X"FE67", X"0100", X"001E", X"0213", X"FF3C", X"FEA6", X"FFA4", X"FF0A", X"FDC9", X"FCB7", X"FE4A", X"FE58", X"005E", X"FED8", X"FFA8", X"0004", X"FEEF", X"007A", X"014C", X"026C", X"04A0", X"0759", X"0689", X"0433", X"04A3", X"FF60", X"FF13", X"0072", X"FF79", X"FC47", X"FB7C", X"0131", X"FE83", X"FF5B", X"FE56", X"FDD0", X"FD21", X"FD69", X"FC1A", X"FBC1", X"FDFB", X"FD1C", X"FDD9", X"00A8", X"FF4A", X"0143", X"038A", X"0355", X"055A", X"06EA", X"0726", X"FFC9", X"015F", X"FCEB", X"0091", X"FF44", X"0005", X"FED5", X"FD4F", X"FD08", X"FF63", X"FE69", X"FD1E", X"FC15", X"FB68", X"FB05", X"FD03", X"FC6E", X"FD7D", X"0070", X"FF8D", X"03DC", X"029D", X"0611", X"072B", X"0741", X"0306", X"04B1", X"01F9", X"0225", X"0112", X"FFEA", X"FF9B", X"00BA", X"0095", X"FE7C", X"01B8", X"021A", X"039B", X"02D1", X"01D9", X"0088", X"0171", X"008B", X"03D2", X"0289", X"0326", X"055F", X"04F1", X"047C", X"0680", X"05BC", X"0756", X"02DE", X"FEAC", X"0137", X"00AD", X"0256", X"0199", X"0263", X"0110", X"014C", X"00CD", X"FE7B", X"FEED", X"FEEA", X"0170", X"03C5", X"06E0", X"069D", X"03F4", X"03D4", X"02E0", X"0479", X"0647", X"05D6", X"0194", X"007E", X"0085", X"0335", X"039F", X"FFAB", X"FDB4", X"FDEB", X"0232", X"007A", X"FF88", X"0034", X"0217", X"FF4E", X"FF44", X"002D", X"FDBF", X"FFE9", X"0160", X"0377", X"05C0", X"03E4", X"034A", X"054F", X"0281", X"056C", X"0A01", X"05E5", X"039D", X"0572", X"0754", X"05B9", X"0530", X"0430", X"0282", X"0037", X"00CD", X"FFF0", X"FDE1", X"0053", X"FEE3"),
        (X"002E", X"FFDE", X"FF87", X"00E8", X"FF67", X"002B", X"009C", X"FEF5", X"FF50", X"FFDE", X"0021", X"0036", X"FFC2", X"FEBF", X"FF68", X"FF39", X"FFB5", X"FF72", X"022F", X"FF75", X"002E", X"FFFF", X"FF07", X"FF0C", X"007D", X"FE8D", X"FFCF", X"FFFB", X"00B2", X"FF7B", X"0052", X"FF67", X"0045", X"FFB3", X"0090", X"0067", X"00D3", X"01D9", X"01A9", X"006A", X"0147", X"FEF0", X"015B", X"FFFC", X"FDF6", X"FDFE", X"013E", X"019F", X"00B6", X"014C", X"FFAA", X"009B", X"0155", X"0086", X"015E", X"FF87", X"00A2", X"FF96", X"FFA3", X"FD7B", X"FEC4", X"0197", X"0158", X"01E7", X"0020", X"FD8D", X"FF5E", X"002F", X"FF6B", X"02FB", X"051A", X"082B", X"0933", X"0967", X"074B", X"07B0", X"06B2", X"04D3", X"03D7", X"0189", X"FDC6", X"FE65", X"FFF6", X"FF77", X"FFF0", X"005C", X"FF88", X"FD35", X"019C", X"0093", X"01EC", X"FDBC", X"FB0B", X"FB8F", X"FAC6", X"F819", X"F824", X"FC54", X"FE46", X"0114", X"0253", X"0344", X"04F3", X"07D5", X"0496", X"0469", X"05A9", X"0107", X"FDD0", X"FC49", X"FD30", X"0019", X"FFEA", X"005C", X"FD76", X"FDD2", X"0018", X"FFF1", X"FD36", X"FCD5", X"FD96", X"FA4B", X"FB6A", X"F7D9", X"F9A2", X"FC11", X"FEC6", X"00BB", X"037F", X"04DC", X"04B6", X"05C2", X"0331", X"0726", X"0436", X"076B", X"0614", X"02E7", X"FF54", X"FF2A", X"01E4", X"FF71", X"00CF", X"FECD", X"028E", X"FF95", X"001E", X"009B", X"FFE2", X"FF08", X"FB5C", X"FA08", X"FBDD", X"FA11", X"FFB5", X"000D", X"00A1", X"0216", X"025B", X"022D", X"053B", X"05BA", X"084C", X"0B17", X"0921", X"0282", X"03C4", X"0132", X"005B", X"00F2", X"FDB5", X"FC37", X"00AE", X"00B2", X"FF48", X"0102", X"FDB0", X"FC15", X"FC16", X"FB09", X"FA2E", X"F9A9", X"F908", X"F949", X"F97A", X"FAC1", X"FCF0", X"FF43", X"00FC", X"0199", X"0498", X"09C9", X"0B35", X"03F8", X"0356", X"FE52", X"FFD5", X"FFE9", X"FA9B", X"FA5C", X"FFAA", X"0139", X"FC80", X"FE8E", X"FB13", X"FBF2", X"FB9A", X"FABC", X"F98E", X"F930", X"F7B2", X"F717", X"F74E", X"F798", X"F991", X"FB4F", X"FCA8", X"FDCF", X"015E", X"0609", X"0915", X"0767", X"02C7", X"FF46", X"FE66", X"FC24", X"FE17", X"FD73", X"FE1B", X"FE0B", X"FD69", X"FCC1", X"F9CD", X"FD3E", X"FB42", X"FB0A", X"F933", X"F8D0", X"F468", X"F310", X"F601", X"F70E", X"FAFF", X"F8F4", X"FC96", X"FB2C", X"FD6F", X"027C", X"0591", X"076E", X"005C", X"0073", X"FF6C", X"FDA3", X"FEEF", X"F948", X"FE9E", X"FB65", X"FBC4", X"FBBC", X"FE44", X"FB48", X"FBC4", X"FBC6", X"FB1E", X"F758", X"F405", X"F618", X"F8E0", X"FAAB", X"FB71", X"FC30", X"FBBE", X"FC7D", X"FC07", X"FC76", X"021F", X"03B5", X"0064", X"FF71", X"0184", X"FFE5", X"FF51", X"FA9E", X"FF6A", X"FC8D", X"FD2D", X"FF76", X"FFCB", X"FE1B", X"FF15", X"FE24", X"FF36", X"FD0A", X"FBE4", X"FFA3", X"FE61", X"FE82", X"FD65", X"FDA9", X"FC3F", X"FBDC", X"FBD3", X"FA50", X"00E7", X"031A", X"0273", X"FE9D", X"01B8", X"FC4E", X"FDFC", X"FFA3", X"009E", X"0127", X"00F3", X"0035", X"01C7", X"024A", X"0234", X"01F7", X"0382", X"038D", X"0543", X"05B3", X"027D", X"FF18", X"FD74", X"FE1B", X"FC6C", X"FAEE", X"FAE1", X"FB14", X"FC0F", X"FE1D", X"FD6C", X"FE45", X"FF9D", X"FCE5", X"0020", X"0145", X"FFF5", X"03C4", X"04F1", X"057F", X"039D", X"03F2", X"0460", X"07FF", X"09C8", X"07A6", X"05B5", X"04B4", X"0215", X"0008", X"FF4F", X"FD86", X"FD1A", X"FE55", X"FD6D", X"008D", X"0015", X"FFF6", X"FE08", X"FDE3", X"0081", X"0028", X"FEE3", X"01AA", X"02BA", X"04C6", X"06D6", X"04A0", X"069E", X"0580", X"073F", X"069A", X"066C", X"04C3", X"0403", X"01F9", X"00CB", X"01CA", X"0129", X"003D", X"FFD8", X"00DD", X"026B", X"05A0", X"0561", X"FFF6", X"FD9B", X"FD48", X"033F", X"008A", X"FD27", X"0162", X"01D8", X"04EE", X"0557", X"04F8", X"0364", X"0461", X"0335", X"049D", X"04BC", X"041D", X"0441", X"02E7", X"0016", X"0314", X"021A", X"0299", X"004F", X"015A", X"0433", X"0417", X"0554", X"FF7B", X"F932", X"FE9C", X"0089", X"019B", X"0405", X"0297", X"0041", X"02B5", X"0310", X"016B", X"03CF", X"01AD", X"FFD7", X"0169", X"030B", X"0476", X"060A", X"033D", X"01E4", X"0221", X"0177", X"02CD", X"01D5", X"0098", X"0258", X"03B4", X"0231", X"FE4F", X"FB77", X"FC3E", X"FF9E", X"0163", X"0097", X"0187", X"FBED", X"0119", X"02F2", X"01AF", X"033F", X"0010", X"FE46", X"FF2A", X"0244", X"05D0", X"07E1", X"03B0", X"012F", X"004A", X"029B", X"03E2", X"0522", X"02D4", X"034E", X"023C", X"FFCF", X"FE3A", X"FD16", X"FBBC", X"005F", X"017D", X"0323", X"FDFE", X"FCBA", X"0104", X"0347", X"020E", X"002D", X"FF34", X"0076", X"008F", X"03A4", X"06DA", X"06CB", X"0429", X"00EF", X"000E", X"0287", X"0415", X"0528", X"02B6", X"0099", X"0159", X"FC9C", X"FD0D", X"FC24", X"FD6D", X"FD2D", X"014E", X"04AF", X"FFBE", X"FEF8", X"FF98", X"0001", X"FFBB", X"FFEA", X"FF32", X"FE52", X"011F", X"055A", X"06A8", X"05AA", X"023F", X"0199", X"0041", X"008F", X"0097", X"0293", X"0084", X"FD6F", X"FDF9", X"FCB4", X"FC8C", X"FDDB", X"0172", X"0052", X"FD6C", X"0392", X"026B", X"FEB8", X"FEC9", X"FF78", X"FE23", X"FE0B", X"008C", X"FEF0", X"01E5", X"030A", X"049F", X"02DA", X"01E8", X"0139", X"FFAE", X"FEC2", X"FE2C", X"004B", X"FEAA", X"FD71", X"FD15", X"FCBB", X"F95E", X"FC51", X"0264", X"FFA5", X"FF06", X"0347", X"01C0", X"FC4D", X"FAE5", X"FE2D", X"FEC4", X"0049", X"0067", X"00E9", X"0296", X"0230", X"0226", X"00F1", X"0197", X"01DE", X"02F6", X"01B3", X"00AF", X"0029", X"FFA2", X"FCE0", X"FB9D", X"FAFB", X"F86A", X"009C", X"00A9", X"0109", X"FFB8", X"FFD5", X"01E3", X"FDE8", X"FC24", X"FE05", X"FDA4", X"FFFC", X"FFD3", X"007E", X"0058", X"FF5A", X"0078", X"01AC", X"0108", X"FFD0", X"045C", X"0242", X"0147", X"0154", X"0138", X"FF5F", X"FD42", X"FC0B", X"FDA9", X"00EA", X"000F", X"01AA", X"00DA", X"0031", X"FF9D", X"0158", X"FD80", X"FBC0", X"FD33", X"FB19", X"FDAD", X"FE39", X"FD78", X"FE60", X"FFAF", X"FF6B", X"0177", X"023E", X"02BB", X"0328", X"034F", X"01BE", X"0066", X"FD6F", X"FDC7", X"FF96", X"FFC4", X"033B", X"0020", X"FE68", X"016A", X"FFD6", X"0008", X"02DC", X"005F", X"FEF1", X"FA37", X"FC7B", X"FF68", X"FE5E", X"FD42", X"FD55", X"FE00", X"FEFB", X"0059", X"FF96", X"0127", X"00FA", X"0019", X"0157", X"FEB1", X"FC8B", X"FACD", X"FEFB", X"02EB", X"0379", X"0055", X"FFEA", X"00CE", X"FF61", X"FDE7", X"FCF4", X"FE16", X"FB85", X"FB7E", X"F8F1", X"FF77", X"FD7E", X"FCD2", X"FD43", X"FC2C", X"FE6F", X"FC1E", X"FB8D", X"FC8D", X"FD87", X"FDB7", X"FE7F", X"FE97", X"FED5", X"FE81", X"FB32", X"0288", X"00F6", X"FFF8", X"0080", X"0063", X"FFEF", X"0025", X"F953", X"F429", X"F809", X"F566", X"F3E2", X"F796", X"F818", X"F8C5", X"F8E2", X"F9B2", X"FA26", X"F8C3", X"F90A", X"F7DF", X"F733", X"F725", X"F65C", X"F723", X"FC49", X"FF3C", X"FD72", X"0013", X"0040", X"FFD2", X"0001", X"FEC6", X"01A9", X"FFFF", X"FD16", X"F92A", X"F683", X"F404", X"F5A8", X"F3A9", X"F2A9", X"F606", X"F5B6", X"F129", X"EE77", X"F46C", X"F2BB", X"F3C6", X"F39D", X"F581", X"F6F1", X"F9A9", X"FA91", X"013A", X"FEA4", X"FF92", X"0025", X"00BC", X"00FD", X"011E", X"FFDD", X"006A", X"FFA0", X"FFD4", X"FBC1", X"FB31", X"FA82", X"FB00", X"FA6E", X"F862", X"F951", X"F988", X"F754", X"F7C3", X"F8AC", X"F9DE", X"F9FD", X"FBAC", X"FC8A", X"FD63", X"FCC7", X"00F1", X"0069", X"005C", X"00CD", X"FFC3"),
        (X"000F", X"FEA0", X"0004", X"0067", X"002E", X"FF9C", X"FF10", X"FFE2", X"00D0", X"FF9D", X"0058", X"FFA8", X"013B", X"0091", X"FF63", X"002B", X"00A3", X"FFC6", X"0034", X"00D2", X"FFC8", X"0031", X"01E8", X"FED1", X"FF82", X"00DE", X"FF3A", X"011F", X"0060", X"FE72", X"FEF6", X"FEE5", X"008D", X"01AE", X"00F9", X"FFEB", X"0241", X"0079", X"008A", X"FFA7", X"0197", X"0065", X"00C6", X"015A", X"0028", X"0008", X"0022", X"0140", X"0236", X"01ED", X"00D1", X"0093", X"FEDD", X"0098", X"00E0", X"FFF6", X"0015", X"00F7", X"FED9", X"FF64", X"FF72", X"0004", X"00D9", X"00FF", X"FF93", X"FDDC", X"0066", X"0051", X"FFF9", X"031A", X"045B", X"0237", X"00E6", X"FED3", X"FE9F", X"FD6F", X"FF8D", X"0189", X"030C", X"FF7E", X"FEEE", X"FF5C", X"0118", X"FFA5", X"FF67", X"008D", X"0012", X"FF17", X"0060", X"0070", X"FE8D", X"FF8D", X"FC9D", X"FE90", X"FE6E", X"FE5E", X"FE07", X"0025", X"0150", X"FF3A", X"FFB5", X"FFAF", X"00CD", X"FFE3", X"FF91", X"0179", X"01B7", X"0136", X"012E", X"FE00", X"000E", X"001E", X"00BC", X"00A3", X"0026", X"FFA7", X"00F4", X"FD1B", X"FCD6", X"F95F", X"FBF2", X"FBE4", X"FEE4", X"FB17", X"FBBB", X"FC9B", X"FB7D", X"FCBD", X"F9FD", X"FB6B", X"FC8E", X"02C7", X"03CA", X"042A", X"028C", X"0351", X"FD2C", X"FC9E", X"FD9C", X"012E", X"006F", X"0042", X"FF1E", X"FF05", X"008D", X"FEAC", X"FDBE", X"FB85", X"FB86", X"FC81", X"FC72", X"F9A6", X"FA62", X"F5EF", X"F98C", X"F8E1", X"F6BE", X"F751", X"F961", X"FAB8", X"FE86", X"FEDA", X"020E", X"02AB", X"00D0", X"FC64", X"0089", X"0213", X"0137", X"010A", X"006B", X"030D", X"0441", X"002A", X"FEEC", X"FDD1", X"FCA4", X"FCDC", X"FCE9", X"FD0E", X"FBE8", X"FA88", X"FBA7", X"FBC0", X"FBF4", X"FA27", X"FBD0", X"FA57", X"FB9C", X"FD18", X"FF51", X"FF51", X"FE9B", X"FD3A", X"FCFE", X"00E3", X"FF64", X"013E", X"0144", X"05F4", X"0375", X"FF6E", X"FF45", X"FD38", X"FBF8", X"FE92", X"FCE3", X"FE1E", X"FEA3", X"FF4D", X"FFA6", X"FE60", X"FE6A", X"FD7C", X"FB19", X"FCEA", X"FC4E", X"FA9C", X"FDA4", X"FDF2", X"FC47", X"FB44", X"FE79", X"014C", X"FFA0", X"03C9", X"00F3", X"02AF", X"0238", X"FF41", X"FEA6", X"FE42", X"FDB3", X"FC40", X"0007", X"0161", X"FF84", X"0091", X"0331", X"0123", X"FF3C", X"009C", X"FE3D", X"FAB9", X"FBC9", X"FBE4", X"FC76", X"FB08", X"F8FF", X"F903", X"F8A6", X"FB50", X"005F", X"04CF", X"0151", X"002B", X"0205", X"FE10", X"FE82", X"FF6D", X"0085", X"001E", X"FFB3", X"01D4", X"026C", X"0248", X"0406", X"05EC", X"026D", X"FEED", X"FFD4", X"FD14", X"FB54", X"FB7A", X"FCB7", X"F97D", X"F9E2", X"F4E6", X"F52D", X"002B", X"016D", X"06C9", X"01C9", X"FF85", X"FF85", X"FD8A", X"FF65", X"012A", X"007E", X"00A0", X"0165", X"003C", X"01C0", X"00AE", X"0541", X"07A0", X"0370", X"0107", X"0137", X"FED8", X"FD1E", X"FD06", X"FC78", X"F9DD", X"F85D", X"F7E4", X"F7B3", X"FFB2", X"003B", X"04FF", X"0272", X"03FD", X"FDBA", X"00A8", X"0241", X"02EF", X"021B", X"020D", X"010D", X"011A", X"FF8F", X"FF56", X"03B7", X"0806", X"04EF", X"02BF", X"02A3", X"00A7", X"FE65", X"FFEB", X"003A", X"FDDD", X"FBCE", X"FABE", X"FA3A", X"0227", X"00F9", X"01BF", X"0481", X"0347", X"0041", X"0208", X"0319", X"05FA", X"00D2", X"024A", X"FF8F", X"00AE", X"FFB0", X"FFDD", X"0344", X"03B7", X"0321", X"016C", X"031A", X"FFF1", X"FF1A", X"00AE", X"032C", X"04C8", X"02CE", X"00F5", X"FBF6", X"023D", X"0043", X"0068", X"02B2", X"0126", X"02AF", X"0416", X"074F", X"0473", X"03C7", X"FFA6", X"FFB2", X"FF06", X"FEA0", X"013F", X"0486", X"020C", X"0221", X"0408", X"0040", X"00FD", X"00B4", X"017E", X"0416", X"0672", X"05BC", X"0246", X"FD63", X"FF4B", X"FFA2", X"01C3", X"0546", X"0355", X"01F0", X"051C", X"0527", X"04D7", X"0382", X"013E", X"0089", X"0108", X"FF23", X"0192", X"0179", X"01E6", X"02C9", X"017A", X"00A6", X"02F2", X"03E6", X"0636", X"064F", X"0717", X"0524", X"0363", X"FD85", X"FD41", X"FFF2", X"FE02", X"0247", X"FE60", X"FFF7", X"0413", X"063D", X"064F", X"0573", X"01C4", X"027E", X"0474", X"0166", X"0067", X"0364", X"0241", X"0337", X"031F", X"02B5", X"0388", X"0538", X"062B", X"0627", X"0709", X"04A5", X"0300", X"FE5E", X"FCF5", X"009D", X"FFBE", X"0070", X"FAC9", X"FDDF", X"00C0", X"05B6", X"0717", X"0790", X"052C", X"04AD", X"05C2", X"038F", X"01D8", X"042E", X"0303", X"034D", X"01C5", X"0150", X"032D", X"043E", X"064F", X"059A", X"039D", X"05FA", X"040F", X"FD3C", X"FDD9", X"00F2", X"018A", X"FE30", X"F973", X"F893", X"FC55", X"01F3", X"05A3", X"06C4", X"0585", X"0779", X"05A5", X"020C", X"04FA", X"06DC", X"050F", X"011A", X"0053", X"FFC9", X"006D", X"01B1", X"0230", X"04B3", X"01AF", X"002D", X"00C0", X"FF4F", X"FB67", X"027C", X"0243", X"012F", X"FACF", X"F768", X"F89A", X"FB46", X"FFED", X"0215", X"03C1", X"04E0", X"0319", X"03B9", X"0563", X"03B4", X"02FD", X"FFBD", X"FF2B", X"00F8", X"FF78", X"004B", X"016F", X"014A", X"FFFC", X"FC31", X"01E0", X"FFF5", X"FE4C", X"013D", X"0188", X"FFF7", X"FC89", X"F91B", X"F697", X"F872", X"FD39", X"FE7D", X"FE9D", X"0012", X"01A7", X"0175", X"FF79", X"0241", X"FF2C", X"0046", X"FEB9", X"FDF4", X"FEC3", X"FF84", X"FF1C", X"FD71", X"FC62", X"FDD2", X"0133", X"FFA5", X"02BD", X"FF2B", X"FF86", X"FFA1", X"FB3E", X"F506", X"F736", X"F9EC", X"FB64", X"FB46", X"FDD2", X"FDD5", X"FFF5", X"005F", X"0182", X"00EC", X"FFB7", X"0089", X"FEA0", X"0096", X"FF02", X"FCB0", X"FAA0", X"F65A", X"F90B", X"018B", X"039B", X"02BF", X"0172", X"002C", X"008D", X"FE0F", X"FBFE", X"FA72", X"FAC3", X"F84D", X"F894", X"FBBA", X"FD04", X"FD08", X"FD76", X"FEE3", X"FDAB", X"0037", X"FE65", X"FF91", X"FFCD", X"FEFF", X"FD63", X"F994", X"F793", X"F28C", X"F863", X"026E", X"0125", X"FF61", X"00A9", X"FFF6", X"00BC", X"FE6C", X"FEF4", X"FF0C", X"0216", X"FC31", X"F9DC", X"FAC8", X"FBCD", X"FBF9", X"F96D", X"F8BB", X"F932", X"FAD1", X"FC5D", X"FC3B", X"FC16", X"FD14", X"FB82", X"F7DF", X"F8DF", X"F4D0", X"F6F7", X"FDAB", X"000A", X"0086", X"FF48", X"FFE5", X"FF97", X"FC37", X"FDE5", X"0092", X"065C", X"032C", X"FFA7", X"FBAF", X"F946", X"FA42", X"F8E8", X"F887", X"FAB5", X"F700", X"F93B", X"F632", X"F9D4", X"FB39", X"FB7A", X"FB03", X"FC1A", X"F91D", X"FA99", X"FD5F", X"FF9F", X"02EA", X"00A7", X"FF3A", X"0059", X"FE1A", X"FED2", X"04E9", X"08F5", X"0552", X"0244", X"FF0A", X"FE3B", X"FF33", X"FA6E", X"F940", X"F928", X"F756", X"F6EA", X"F826", X"FD93", X"FF38", X"FF52", X"FFBA", X"045C", X"FF4D", X"0111", X"FC70", X"01D0", X"FFCA", X"FEDA", X"00EC", X"0038", X"FF0D", X"030D", X"0286", X"05EE", X"03B7", X"0689", X"0712", X"03BB", X"0340", X"0220", X"0296", X"FFF0", X"FF1D", X"FDA6", X"FE57", X"FFE6", X"FE9C", X"FF5A", X"0203", X"03A3", X"00BB", X"FE7C", X"FEF4", X"0174", X"010B", X"00C6", X"00C7", X"FFB1", X"0012", X"FFB3", X"00D2", X"03C3", X"05F2", X"06AA", X"0705", X"07A9", X"0871", X"0512", X"04D5", X"0606", X"0C5D", X"0869", X"07CB", X"05DB", X"01D8", X"01B6", X"0068", X"FFB1", X"0028", X"FF80", X"0047", X"007E", X"00AC", X"FF9F", X"0155", X"00B5", X"FF47", X"00B5", X"00BA", X"008E", X"022C", X"01D9", X"0143", X"0303", X"03CA", X"01EF", X"02DD", X"04B8", X"067C", X"06C5", X"04AE", X"03A4", X"04D9", X"037E", X"0274", X"031D", X"0199", X"00A9", X"FF70", X"004F", X"FFB1", X"0017"),
        (X"FF74", X"FFEF", X"FE6D", X"FF74", X"FFCE", X"003D", X"0022", X"0057", X"0037", X"FF96", X"0109", X"0114", X"FF0B", X"FD00", X"000B", X"FF5E", X"0186", X"FFE1", X"FFB7", X"FF80", X"FFA4", X"FFB8", X"FF9D", X"010B", X"FFA9", X"00DB", X"01C2", X"FF55", X"008A", X"012D", X"006A", X"007E", X"0015", X"005A", X"FDCD", X"FDDA", X"FCBF", X"FA99", X"FA65", X"FA14", X"F997", X"F9C2", X"001E", X"FE5B", X"FB07", X"F9AF", X"FBC3", X"FC69", X"FB19", X"FAD2", X"FC68", X"FE88", X"FFF8", X"FFDE", X"00BF", X"0014", X"00DD", X"0033", X"FEFF", X"FC40", X"FE03", X"FF35", X"FAF6", X"FA1A", X"FA09", X"F71A", X"F6C0", X"F3C3", X"F4CA", X"F879", X"F691", X"F7F1", X"F81E", X"FB22", X"F753", X"F82E", X"FA64", X"FAB5", X"F9CC", X"F8B2", X"FBB1", X"FDF4", X"0003", X"FF24", X"0088", X"0020", X"01AA", X"FD3B", X"FD47", X"FB82", X"FA20", X"F4FA", X"F6B1", X"FA01", X"F5D0", X"F7A0", X"F5F0", X"F311", X"F357", X"F7A7", X"F88A", X"F687", X"FA35", X"FB00", X"FA02", X"FD64", X"FD30", X"FAD5", X"FB30", X"FF0C", X"FD2F", X"004A", X"00F7", X"FF6A", X"036D", X"01F2", X"015B", X"00BB", X"FCCD", X"FAF1", X"FC2B", X"FC86", X"FA98", X"FA37", X"FB22", X"FD01", X"FBCD", X"FCBB", X"FECA", X"FFE3", X"FCD5", X"FDB8", X"FCD8", X"FE56", X"FDD4", X"0046", X"FFE5", X"FE1F", X"0202", X"FD24", X"FECE", X"0130", X"FE04", X"FF67", X"FFFF", X"0269", X"FE27", X"FCC8", X"FD10", X"FC26", X"FA5B", X"F9B5", X"FCD9", X"FA7D", X"FC0C", X"FC0F", X"FC97", X"FB6F", X"FB29", X"FE3E", X"0044", X"015F", X"018F", X"0232", X"0332", X"0164", X"0035", X"FDB7", X"005C", X"FF7A", X"FF9C", X"0025", X"007A", X"0271", X"FDEE", X"FDA2", X"FBDB", X"FCC3", X"FC9E", X"FAD9", X"FB88", X"FA87", X"FC5F", X"FCBD", X"FB3E", X"FE73", X"FEAA", X"0332", X"02F4", X"00E5", X"0462", X"04BD", X"0426", X"05D8", X"088F", X"022A", X"0061", X"0170", X"FFBD", X"0332", X"FFFE", X"00CA", X"FD79", X"FF67", X"FDBB", X"FBCD", X"FD70", X"FEF7", X"FDF0", X"0074", X"FEC5", X"FEC3", X"FF98", X"00A4", X"041D", X"04DF", X"03CE", X"03E3", X"051E", X"04CF", X"0311", X"031A", X"04AB", X"02B3", X"FD6C", X"00AA", X"0143", X"FFA6", X"003B", X"0345", X"014D", X"FFE5", X"FE78", X"FF72", X"FF73", X"022E", X"0391", X"03A4", X"01FB", X"01AE", X"0369", X"0357", X"0416", X"02BC", X"03AE", X"039E", X"01D3", X"0549", X"0704", X"0B31", X"06BB", X"035F", X"FF94", X"00CF", X"FDEF", X"FFC5", X"FF99", X"0146", X"FFFE", X"FEFE", X"0080", X"00E1", X"01B8", X"04AC", X"0518", X"059C", X"01A8", X"0134", X"0139", X"031F", X"03DE", X"0231", X"0147", X"01CB", X"00C9", X"051C", X"0742", X"0B62", X"05E2", X"02BE", X"FF48", X"012A", X"FD34", X"0022", X"04DC", X"0092", X"02C1", X"026D", X"02A6", X"065C", X"060C", X"0728", X"07FD", X"025A", X"038B", X"025D", X"025D", X"010B", X"035C", X"0281", X"FFAF", X"0247", X"01DF", X"FF4D", X"04F9", X"0953", X"0721", X"0335", X"0263", X"018D", X"0200", X"0174", X"05E2", X"06AC", X"0779", X"09C0", X"06E7", X"068F", X"05EC", X"0640", X"0473", X"018E", X"0209", X"0346", X"03A8", X"00CF", X"00BC", X"FF4B", X"FD7D", X"FDF4", X"0087", X"FD08", X"FF7D", X"0422", X"06C2", X"03D7", X"00E6", X"01AE", X"02D8", X"0485", X"061A", X"0938", X"0929", X"0AAE", X"06A4", X"063B", X"0425", X"01BD", X"FDDB", X"FF16", X"02D4", X"013B", X"00D4", X"0032", X"0033", X"FE71", X"FEB7", X"FF74", X"FEBF", X"FC8C", X"FCBB", X"FF4C", X"0157", X"FEA8", X"FFA8", X"024E", X"0417", X"020F", X"04FF", X"060F", X"0541", X"068C", X"04A4", X"0329", X"FE80", X"FB27", X"FA81", X"FEEF", X"0257", X"02BE", X"007F", X"0128", X"FF31", X"FDDD", X"000F", X"FFBD", X"FD9D", X"F807", X"F685", X"FB56", X"FA3D", X"FAE1", X"0340", X"00F1", X"0428", X"FEDE", X"04E4", X"0297", X"01C5", X"00D8", X"030B", X"00C4", X"FADB", X"F6C9", X"FAED", X"01A5", X"03C2", X"0360", X"0227", X"03F2", X"FF48", X"FF4E", X"FDAE", X"FC5E", X"FCC5", X"F891", X"F6FF", X"F95B", X"F8B9", X"FD14", X"0254", X"005B", X"0102", X"0015", X"FE12", X"FD03", X"FE39", X"FD9A", X"0124", X"FEDA", X"FA8B", X"FBF8", X"01E8", X"0606", X"057E", X"0536", X"0245", X"02C3", X"FF32", X"FAC5", X"FB4B", X"FB0C", X"FBA2", X"F8AD", X"F6DE", X"F505", X"F8CB", X"FE84", X"0086", X"FFD7", X"FCBB", X"FBEA", X"FA73", X"FA5E", X"FE2F", X"FDC3", X"0043", X"FED6", X"FF8D", X"0222", X"067A", X"0639", X"0527", X"04EC", X"0397", X"0143", X"FC24", X"FB5F", X"FC05", X"FDA2", X"FB3D", X"FB1A", X"F721", X"F448", X"F95C", X"FEEE", X"FFC4", X"00A9", X"FDFE", X"F96F", X"F888", X"FB37", X"FA7D", X"FCA9", X"FE2A", X"0115", X"01B4", X"03EB", X"05D9", X"063D", X"0623", X"03A7", X"02FF", X"FD2D", X"FD32", X"FBA2", X"FC8A", X"FC81", X"FB9A", X"FAB4", X"F77F", X"F6CF", X"FBE3", X"FE0C", X"0042", X"004E", X"FD57", X"F7BA", X"F72F", X"F8FA", X"FA60", X"FA65", X"FB1F", X"FF6E", X"FE5B", X"FF4D", X"00F4", X"0434", X"0456", X"0084", X"FC6E", X"FCB8", X"FC3C", X"FD3B", X"FDC9", X"FE0E", X"FA5E", X"F656", X"F7F9", X"F768", X"FEFF", X"005E", X"FF7E", X"FED1", X"FF95", X"F60F", X"F63A", X"F9A5", X"FA88", X"FB79", X"FA88", X"FA9C", X"F8B6", X"F93C", X"FC56", X"FE73", X"0131", X"FD2C", X"FDF3", X"FF74", X"FDF9", X"FCFB", X"FCB4", X"FE6B", X"FCA4", X"FA90", X"FA65", X"F8E8", X"00AB", X"0270", X"026C", X"FD2B", X"FAF3", X"F593", X"F3D3", X"FA52", X"F9F1", X"FB2A", X"FB06", X"FA28", X"F960", X"F8EA", X"F903", X"FAA2", X"FC5E", X"FC4D", X"FE8F", X"FF8A", X"FF34", X"FF0D", X"FE89", X"FD2D", X"FE12", X"FC15", X"FAFE", X"FB7A", X"0057", X"00B7", X"00FE", X"FF89", X"FACB", X"F77A", X"F93E", X"FB6D", X"FCD8", X"FCC0", X"FAB5", X"FA6B", X"FAB1", X"FA4F", X"FA34", X"FAC3", X"FC40", X"FF07", X"FD22", X"FF5B", X"FD7A", X"FC6C", X"FE10", X"01B6", X"FFC4", X"FC9A", X"FD27", X"FF27", X"FB6A", X"FFA0", X"00C2", X"FFFA", X"FB3E", X"F7B7", X"FDAF", X"FE73", X"FCAF", X"FFA9", X"FD3C", X"FDC6", X"FD38", X"FDCD", X"FD39", X"FC7F", X"FFC6", X"FDD1", X"FF80", X"00D2", X"FE7B", X"FB35", X"FC5A", X"0031", X"FD0D", X"FDBA", X"FF24", X"FFF9", X"026B", X"00A3", X"FDCF", X"00C2", X"FD73", X"F949", X"FB46", X"FFD5", X"00B7", X"FE64", X"0033", X"FFF9", X"FFEE", X"00EA", X"00C8", X"0122", X"0227", X"00F1", X"00E3", X"FF04", X"FD4F", X"FDBC", X"FF31", X"0030", X"FE8A", X"FFC7", X"FDCB", X"FBA8", X"022E", X"FF3E", X"0016", X"0086", X"FEEA", X"FA08", X"F9AA", X"0027", X"FF15", X"FFB0", X"FF89", X"FFD6", X"FF11", X"FF73", X"FF89", X"FED7", X"FF35", X"FF95", X"FD2F", X"00D9", X"FEEF", X"0044", X"FD90", X"FDCA", X"FF03", X"00EB", X"FBD1", X"FCCF", X"FDC2", X"FF91", X"FF70", X"FF39", X"FCFF", X"0185", X"0259", X"01D7", X"0214", X"0569", X"047C", X"0412", X"02D8", X"021E", X"0323", X"021E", X"024F", X"0479", X"0190", X"0080", X"FD53", X"FAB9", X"FDB6", X"0060", X"FFEA", X"02D1", X"FF01", X"FF7C", X"FFB2", X"FF1F", X"01D2", X"0134", X"0053", X"FEA9", X"FDB6", X"00FC", X"0259", X"05EA", X"0922", X"064B", X"079A", X"077F", X"044A", X"0375", X"04F0", X"06CB", X"04CE", X"0546", X"044F", X"FFD8", X"FFB9", X"023A", X"00C2", X"0113", X"FF38", X"FEB9", X"0077", X"FF0D", X"01D8", X"005E", X"FE52", X"FEB1", X"FF8E", X"00EC", X"0126", X"0064", X"019D", X"0131", X"01DE", X"00BA", X"00AF", X"028A", X"020F", X"0177", X"0281", X"0150", X"018A", X"0326", X"034A", X"03B4", X"013F", X"0202", X"FFD0", X"0030", X"FF85", X"02D3"),
        (X"FF80", X"FF93", X"FF4E", X"FEDB", X"0042", X"0043", X"00C7", X"FEF5", X"FF5E", X"0032", X"00A3", X"007B", X"0002", X"01B2", X"00A0", X"FF9C", X"FF66", X"FFB5", X"00CC", X"004E", X"FF74", X"0086", X"0154", X"FF8A", X"012F", X"FE93", X"00B3", X"FFC3", X"FF23", X"0072", X"0003", X"FFF6", X"004B", X"001E", X"042A", X"04E6", X"0476", X"0563", X"060E", X"03EB", X"05F6", X"052B", X"FF75", X"00DC", X"0000", X"05CC", X"060E", X"0613", X"064C", X"0573", X"03DD", X"03F3", X"FEF0", X"FF4F", X"0093", X"00DD", X"FE2D", X"FFA8", X"00EF", X"FFFD", X"01D7", X"00A3", X"036F", X"057E", X"0521", X"0750", X"0812", X"093E", X"0888", X"0ADB", X"09C8", X"0590", X"0406", X"04EC", X"0712", X"0A6F", X"0895", X"08B3", X"07FE", X"05C3", X"FE7D", X"FF05", X"FFF2", X"0138", X"FEF9", X"FE9D", X"0039", X"0301", X"0243", X"03B2", X"05E8", X"0525", X"055D", X"0820", X"0630", X"08F5", X"081C", X"0A15", X"078A", X"06F5", X"05B3", X"059C", X"063E", X"0544", X"057C", X"038C", X"0409", X"052D", X"00E4", X"FF38", X"FFD4", X"FF64", X"000C", X"00BD", X"0149", X"0311", X"0444", X"050D", X"0460", X"051B", X"04CD", X"03E3", X"03D1", X"0159", X"0026", X"FFCE", X"FE0D", X"FFA0", X"0178", X"0103", X"027F", X"061A", X"0783", X"045F", X"06D7", X"0625", X"01AD", X"FF29", X"FF57", X"028A", X"FF2D", X"FFAB", X"02E7", X"00BB", X"049A", X"03D5", X"03FD", X"0299", X"0186", X"00B6", X"0363", X"004F", X"FF3C", X"FEB0", X"FDC6", X"00EB", X"012B", X"FF93", X"0126", X"0384", X"0636", X"054B", X"058F", X"0B11", X"0A27", X"0481", X"02CF", X"0220", X"014D", X"0115", X"FE7B", X"036A", X"072F", X"02DA", X"0278", X"004F", X"002D", X"FF61", X"0044", X"0035", X"FFA3", X"FFA7", X"0005", X"FEAE", X"FD68", X"FCEC", X"FDF2", X"FFDB", X"FF3E", X"0159", X"0373", X"06F9", X"0AD2", X"08B3", X"0566", X"028B", X"FF03", X"01DE", X"FD75", X"FF97", X"0505", X"0173", X"007D", X"FEFE", X"FE0A", X"FD71", X"FD97", X"FBAD", X"FDD4", X"FB25", X"FDA6", X"FD46", X"FCD8", X"FB81", X"FBC0", X"FC49", X"FB59", X"FBDA", X"FC3E", X"FEEC", X"048B", X"06D0", X"072C", X"0158", X"0160", X"FF95", X"FD12", X"FF04", X"02D0", X"FF3C", X"FCAB", X"FCF5", X"FE1E", X"FA80", X"FBF0", X"FA47", X"F9D6", X"FA0B", X"FBD2", X"FC0B", X"F98D", X"FB2D", X"F7E7", X"F9A4", X"F9FB", X"F92C", X"F871", X"F661", X"FBBC", X"01A0", X"01E9", X"FC2B", X"FFAC", X"FE6D", X"F9EE", X"FDBC", X"023A", X"FA97", X"FBC9", X"FD49", X"FCA5", X"FBD9", X"F9FF", X"F8AA", X"F8DE", X"F89E", X"FC30", X"FD4D", X"FCDA", X"FB25", X"F905", X"F8C3", X"F9DC", X"F98A", X"F924", X"F803", X"FBF5", X"0592", X"0202", X"FF7D", X"00B5", X"010C", X"FAB6", X"FDED", X"FE7D", X"FAD2", X"FC4E", X"FBC8", X"FA00", X"F767", X"FB31", X"FA5C", X"FACC", X"FDD6", X"009F", X"01C5", X"0093", X"FDEE", X"FAB3", X"FC47", X"FDBB", X"FBBF", X"FF46", X"FF5E", X"01A6", X"040C", X"FEE4", X"FE16", X"0035", X"FE34", X"FF26", X"FE6C", X"FE49", X"FD2F", X"FF9D", X"FD26", X"FCDD", X"FCC8", X"FBDD", X"FEBE", X"0313", X"0483", X"0434", X"039A", X"0342", X"FEFA", X"FD35", X"FD70", X"FD4B", X"FEDE", X"00BD", X"031F", X"01C1", X"00DA", X"FCA8", X"FEC2", X"FFBA", X"FE1B", X"FC15", X"FB12", X"FE5F", X"FEBB", X"01F0", X"0193", X"0088", X"016C", X"026A", X"0430", X"04C5", X"0294", X"04C4", X"039E", X"0301", X"FF9F", X"FE9A", X"FD70", X"FE6E", X"FFF8", X"FFBB", X"031F", X"01F3", X"00BD", X"F881", X"FD97", X"01D4", X"FE6D", X"FCC4", X"FD8C", X"FFAD", X"0109", X"0508", X"02C1", X"040F", X"0311", X"034D", X"0137", X"0288", X"0309", X"04C8", X"0355", X"03C4", X"FEFA", X"FCEE", X"FF09", X"FE61", X"0055", X"0255", X"055B", X"031E", X"FCC9", X"F82D", X"FD4C", X"FF0F", X"FFBB", X"002C", X"FFB8", X"FBAC", X"01DC", X"025F", X"00F7", X"0152", X"03FC", X"0119", X"FEBD", X"0060", X"02EE", X"01A5", X"00F4", X"0208", X"FD8B", X"FE3C", X"FFFA", X"FEFC", X"0216", X"0528", X"0467", X"01F0", X"FEB6", X"F8A1", X"FD0E", X"006B", X"006A", X"04D5", X"FCBA", X"F8F5", X"FF41", X"006F", X"FF37", X"FD5D", X"FE8D", X"FD73", X"FE3F", X"0055", X"042F", X"0316", X"0181", X"FDC4", X"FC04", X"00C4", X"03D0", X"019A", X"0386", X"035D", X"02D2", X"0057", X"FF4E", X"F76D", X"FCC1", X"FF24", X"023B", X"0504", X"FE91", X"FBC1", X"FC72", X"FBE4", X"FC3F", X"F966", X"FB97", X"FCBD", X"FCDA", X"FD40", X"0308", X"036B", X"FC6D", X"FC12", X"F94B", X"FF34", X"03F2", X"0303", X"0077", X"037A", X"028C", X"005A", X"FB7F", X"F7AA", X"FBCC", X"003B", X"01C2", X"04CF", X"FF58", X"FA66", X"FC3F", X"FB39", X"FBB4", X"FBA9", X"FB85", X"FDF4", X"FCF8", X"FC34", X"000A", X"FF4B", X"FC11", X"FB9D", X"FD38", X"00CA", X"03BB", X"0252", X"00C2", X"006A", X"0208", X"FE5C", X"FC0D", X"FA3A", X"FDE3", X"FEA2", X"0019", X"05B5", X"05D5", X"FC93", X"FAC1", X"FBB6", X"FD3A", X"0007", X"015C", X"00CF", X"FFCA", X"0203", X"0152", X"FF4F", X"FDDE", X"0137", X"02DA", X"01AB", X"00FB", X"0194", X"0230", X"0258", X"0151", X"FE52", X"FE2D", X"FAE0", X"0025", X"00B8", X"FDD2", X"075F", X"07FE", X"FE5B", X"FA42", X"FEF0", X"FE5F", X"00FC", X"0320", X"0595", X"0447", X"03FF", X"0567", X"0239", X"0331", X"03E2", X"0505", X"024C", X"FFE0", X"011F", X"011F", X"0106", X"FF9F", X"FE2E", X"FD6A", X"FE02", X"00C9", X"0020", X"FF34", X"04B9", X"082B", X"FFF4", X"FD44", X"01CC", X"00D9", X"0193", X"043E", X"05D1", X"0675", X"03C7", X"03E6", X"060B", X"02C3", X"0501", X"02F1", X"03E7", X"0241", X"03AD", X"0133", X"FE60", X"FD92", X"FCA0", X"FA74", X"029F", X"0176", X"0121", X"00E7", X"037C", X"0467", X"0276", X"0125", X"023F", X"0343", X"023A", X"0266", X"0479", X"0262", X"028C", X"0410", X"05D5", X"05EC", X"042D", X"04DF", X"0599", X"046A", X"035D", X"FEE2", X"F967", X"F7A2", X"FB0D", X"FC3B", X"0027", X"00B8", X"00F0", X"01A4", X"0325", X"024D", X"00B7", X"0569", X"0133", X"0046", X"0085", X"FFCE", X"FEFC", X"FF70", X"FE64", X"FDED", X"00A9", X"031C", X"03FA", X"041D", X"0468", X"02A5", X"00FD", X"F94E", X"F4FA", X"F44E", X"F6C0", X"FDC5", X"032F", X"FFD7", X"020D", X"0280", X"038C", X"01EB", X"0528", X"0678", X"048B", X"01A5", X"007D", X"0319", X"00B2", X"FDA8", X"FC49", X"FD77", X"FCEB", X"0167", X"FEEE", X"0056", X"0004", X"FE77", X"FBCD", X"F8E8", X"F8B7", X"F58A", X"FC9A", X"FEEB", X"043E", X"0082", X"0171", X"0038", X"0047", X"0247", X"02E4", X"04C9", X"027F", X"00E9", X"00A6", X"02EE", X"00B3", X"005D", X"009A", X"FFDF", X"FEB0", X"FBC6", X"FAA9", X"FC62", X"FA0B", X"FBF7", X"F7A1", X"F8A1", X"F9AF", X"F8BF", X"FB6E", X"015E", X"02CC", X"0118", X"FFE9", X"FF52", X"0212", X"0076", X"FDF1", X"FD2C", X"FD63", X"FC44", X"FD0A", X"FCDA", X"F806", X"F8D5", X"FCBA", X"FAEB", X"F9B8", X"F712", X"F6AE", X"F770", X"F53E", X"F71A", X"F8E0", X"FC25", X"FCE2", X"FB7C", X"FCDD", X"FE73", X"006C", X"FF73", X"FEF6", X"FF8F", X"FF93", X"FF43", X"FD89", X"FDA2", X"FD51", X"FD25", X"FB63", X"FB6A", X"FA0D", X"FB12", X"F893", X"F92B", X"F7C9", X"FA6E", X"FA8A", X"F729", X"F779", X"F979", X"FE9C", X"FF3B", X"FFF4", X"FFC2", X"0063", X"01D7", X"0079", X"FECA", X"FE99", X"0136", X"FFFE", X"FF1E", X"FE03", X"FF58", X"FFA1", X"FF06", X"FEAC", X"FDD8", X"FDA8", X"FE6A", X"FE1B", X"FB84", X"FCC0", X"FC9C", X"FF1E", X"FDEA", X"FBFA", X"FDC1", X"FFDA", X"FF90", X"005B", X"FF13", X"FF98", X"FF66", X"002E", X"0125"),
        (X"FF4B", X"FF2E", X"FF3E", X"FF9E", X"FEC6", X"0011", X"0081", X"FFE5", X"013A", X"0048", X"FFF4", X"0116", X"FDF8", X"FE1B", X"0047", X"008E", X"FF29", X"FFC8", X"FF71", X"FFFC", X"0134", X"00A9", X"FD8B", X"FEC6", X"001C", X"0073", X"0014", X"0110", X"00C5", X"FE91", X"FFD1", X"012B", X"FF50", X"FFCD", X"003B", X"0019", X"0066", X"FE94", X"FC78", X"FDB5", X"FD06", X"FC13", X"FEF8", X"FC07", X"FD6A", X"FCF5", X"FA2E", X"FD1D", X"FBC5", X"FF79", X"FD3E", X"FD84", X"FFAF", X"FF07", X"FFBB", X"FFDB", X"015A", X"0079", X"015C", X"FF52", X"FD18", X"0009", X"FF10", X"FF5D", X"FF67", X"0292", X"01A9", X"FF4C", X"0128", X"FD72", X"FEFF", X"FEB7", X"FD98", X"FE48", X"FB18", X"FA76", X"FC81", X"FB26", X"F8FA", X"F928", X"FF34", X"01B7", X"FFA8", X"FE93", X"0065", X"FFF4", X"0084", X"FE14", X"FE1E", X"0254", X"0319", X"038C", X"07D1", X"097C", X"08DE", X"0BA0", X"0591", X"0342", X"029E", X"0044", X"00A2", X"FF69", X"FC2F", X"FD6F", X"FCBF", X"F844", X"F8BB", X"F958", X"FCBF", X"02E9", X"FD7B", X"006B", X"0115", X"FED4", X"0170", X"032B", X"0573", X"0671", X"08CE", X"097C", X"0965", X"06E2", X"0478", X"049A", X"04A3", X"0490", X"01DD", X"FDF3", X"FBFD", X"FC9A", X"FC9F", X"FE41", X"FD42", X"FA3A", X"FC4F", X"F8B6", X"FE25", X"FEF6", X"FB95", X"FC5F", X"00B9", X"0014", X"00E1", X"04DE", X"075C", X"091D", X"0D09", X"0BB9", X"07EC", X"030B", X"01B2", X"015D", X"01F9", X"029C", X"0126", X"01CF", X"001E", X"FDE4", X"FE18", X"FEA2", X"FE9B", X"FC36", X"FE09", X"FC21", X"FBAA", X"FE2D", X"FC7B", X"FD5A", X"FF7D", X"0013", X"0049", X"0614", X"079B", X"0B59", X"0E58", X"090A", X"0654", X"0199", X"0285", X"FDD7", X"0017", X"0011", X"007A", X"FFFB", X"0012", X"FFBE", X"FD82", X"FB84", X"FBB6", X"FF11", X"FEE4", X"FC30", X"FCB0", X"FA8F", X"FBD0", X"FDE5", X"FE14", X"00F0", X"00D3", X"06FE", X"0998", X"0BEA", X"0C79", X"0696", X"02EE", X"005A", X"FF60", X"FE08", X"FE24", X"FF23", X"FF5B", X"FF68", X"00A5", X"FE8B", X"FBCC", X"FD42", X"FA8B", X"FA96", X"FAD2", X"F942", X"FA66", X"F7FD", X"FE4D", X"FD1F", X"00F1", X"001C", X"040D", X"08E1", X"0ABA", X"0ADE", X"08B6", X"03F0", X"01D9", X"FE72", X"FF7D", X"FD33", X"FEC2", X"0128", X"FF8C", X"0208", X"01CD", X"FEB0", X"FE20", X"FA25", X"F902", X"F9D6", X"F9A5", X"F882", X"F61E", X"F67A", X"FA31", X"FE5B", X"014D", X"00A5", X"038E", X"071E", X"072E", X"070E", X"0799", X"03CB", X"FF1F", X"FD79", X"FD3A", X"FB37", X"FE60", X"FDFF", X"01F3", X"0405", X"049C", X"0467", X"051C", X"03E3", X"0037", X"FCA2", X"FB29", X"F9B9", X"F4C5", X"F2AC", X"F815", X"019D", X"FFD3", X"026D", X"0339", X"06F3", X"055E", X"04D8", X"04C0", X"00BC", X"FD27", X"FD9C", X"FD21", X"FC92", X"FD76", X"FEC1", X"FF8D", X"03A9", X"086F", X"0AD4", X"0DBF", X"0F51", X"0CD9", X"07A6", X"05EA", X"0083", X"FB6D", X"F68E", X"F815", X"0072", X"012D", X"01EE", X"0395", X"0857", X"0259", X"015E", X"0016", X"FF80", X"FE68", X"FFD4", X"FF8B", X"0283", X"FF2C", X"FDC6", X"FF09", X"0335", X"0722", X"0A6D", X"0F35", X"15C1", X"188E", X"1544", X"1214", X"0DA1", X"07A6", X"FA1F", X"F8EB", X"00C4", X"FF9E", X"04C3", X"0559", X"01D8", X"01E1", X"00BA", X"FE68", X"FF9C", X"00D6", X"0307", X"025B", X"01A4", X"01AE", X"00B1", X"FDF9", X"0308", X"06C6", X"053D", X"0510", X"0A93", X"1463", X"17C2", X"16F4", X"142C", X"1161", X"0426", X"0036", X"FF73", X"FDE1", X"0008", X"023B", X"FEE2", X"FE74", X"FE3E", X"003B", X"003D", X"0151", X"000B", X"0327", X"0242", X"01B7", X"FD3A", X"FD91", X"0260", X"046F", X"0110", X"FF60", X"FD91", X"032A", X"1150", X"1531", X"143B", X"105D", X"084F", X"FDB0", X"FF9F", X"FE04", X"0149", X"0208", X"03B6", X"00DD", X"0218", X"FF4D", X"015B", X"0020", X"FE22", X"FF5F", X"0179", X"0067", X"FFF8", X"FEB8", X"01E9", X"0324", X"0277", X"FE0C", X"FBBB", X"FAE3", X"052D", X"0FFC", X"1208", X"0F5A", X"0658", X"01D0", X"FEEE", X"FE4A", X"02B9", X"02AD", X"0365", X"04E0", X"033B", X"0244", X"0427", X"FF96", X"FE12", X"FF84", X"006B", X"FE4E", X"FF30", X"01A6", X"031D", X"0203", X"0181", X"FE73", X"FDEE", X"FCAF", X"002A", X"0864", X"0E2A", X"0B69", X"058D", X"03E0", X"0466", X"0254", X"004B", X"0340", X"01BC", X"0257", X"0401", X"04AE", X"04A8", X"0256", X"01C8", X"0025", X"FE6C", X"FF81", X"0068", X"FF93", X"03D7", X"0128", X"0074", X"0018", X"007B", X"0016", X"00F1", X"03B9", X"09E8", X"0A46", X"06C7", X"0283", X"049D", X"00AA", X"00E3", X"020F", X"FEC7", X"FF32", X"0010", X"003C", X"03B2", X"02A3", X"01E3", X"012C", X"FDED", X"FFE0", X"0169", X"00AB", X"00FE", X"0296", X"FFEF", X"FF17", X"FE54", X"FE17", X"FFB2", X"01DC", X"079A", X"07DE", X"0A7E", X"02C3", X"0318", X"FFCE", X"0334", X"01F4", X"0044", X"FC83", X"FE98", X"FDE7", X"0039", X"014A", X"0061", X"010A", X"0065", X"FE1C", X"005F", X"FF90", X"FFD6", X"FF7D", X"FE57", X"0001", X"003B", X"FE85", X"FF8A", X"0145", X"0417", X"065E", X"073C", X"047E", X"0218", X"FF5F", X"0385", X"FCF3", X"015F", X"FE52", X"00A8", X"0154", X"00A3", X"FDDA", X"FD9D", X"0057", X"FDF8", X"FE59", X"FF89", X"005A", X"008F", X"00ED", X"0176", X"009A", X"0176", X"0025", X"FE9D", X"FE5E", X"0220", X"0056", X"04EA", X"0413", X"0106", X"01E8", X"02F7", X"FEC5", X"00F9", X"FFF4", X"FE90", X"00E4", X"000E", X"FD45", X"FDB6", X"FC72", X"FC36", X"FD84", X"0122", X"0056", X"FE8E", X"0069", X"FD90", X"FEB1", X"FE28", X"FDAE", X"FDC9", X"FC7E", X"025C", X"FF09", X"0654", X"0092", X"00CF", X"FF7A", X"02C1", X"0752", X"01A3", X"FC66", X"0057", X"000D", X"FEBC", X"FF0D", X"FDE3", X"FEDC", X"FEC5", X"FF23", X"FDC4", X"FE9D", X"FE30", X"FEA6", X"FE6B", X"FE43", X"FE38", X"FBEF", X"FB00", X"FC8B", X"009D", X"01F0", X"02C3", X"00F8", X"FED3", X"0098", X"FF3D", X"05C2", X"00CF", X"FB48", X"FE0E", X"0123", X"01C0", X"FF64", X"FF7E", X"0013", X"FF53", X"FF67", X"0047", X"FF53", X"FDFF", X"FF0B", X"FEB9", X"FE42", X"FBFE", X"FB31", X"FC79", X"FF4A", X"FEF5", X"00F2", X"FFCF", X"FB12", X"0135", X"FFC7", X"FEF3", X"023C", X"FFDF", X"FE7E", X"FB97", X"FE3F", X"0184", X"FFB2", X"FF25", X"FF3D", X"028D", X"00EE", X"0097", X"0124", X"FF6C", X"FF06", X"FFBE", X"FDF7", X"FDFF", X"FC53", X"0068", X"FEA3", X"FE20", X"FF56", X"FF3A", X"FDF1", X"0073", X"0097", X"FFE4", X"0217", X"FF28", X"0393", X"02EC", X"FD53", X"FFBD", X"FF26", X"FF25", X"0180", X"0106", X"FFEE", X"008B", X"0121", X"00D7", X"0253", X"0037", X"FFCA", X"FEA5", X"FE38", X"0032", X"FDFA", X"FF4F", X"FD06", X"FE7B", X"FE92", X"FF36", X"0089", X"008E", X"00D5", X"FD2D", X"0109", X"04D7", X"013D", X"FF98", X"FFB0", X"FF9B", X"0089", X"FDC7", X"FCC2", X"FD45", X"008B", X"FE8E", X"FDD6", X"FE67", X"FF29", X"01F6", X"0109", X"FE9B", X"FD98", X"FD2E", X"FC5A", X"FEF2", X"FE5F", X"FFAE", X"002E", X"0084", X"FFB3", X"0062", X"0214", X"0149", X"05A5", X"0770", X"0582", X"01DB", X"FFFC", X"FF19", X"00DE", X"019B", X"017A", X"000F", X"FFEA", X"01CB", X"0443", X"01DA", X"FFAA", X"FECA", X"FD7C", X"FEC4", X"0008", X"002A", X"001D", X"FFA2", X"FFE8", X"0033", X"FF7C", X"005D", X"01C6", X"00A2", X"00E1", X"FF12", X"015F", X"006C", X"FF55", X"FDE5", X"000A", X"01B9", X"0345", X"03DD", X"0337", X"0136", X"0417", X"03D5", X"00D4", X"008E", X"01F9", X"0043", X"FF94", X"FED4", X"019A", X"FFDE"),
        (X"00E9", X"006A", X"0081", X"006D", X"FDAA", X"0023", X"FF5B", X"0081", X"FFE5", X"0044", X"0037", X"003F", X"0008", X"0124", X"FF2C", X"007E", X"00B2", X"FF86", X"FFF9", X"0036", X"FF34", X"006D", X"FF99", X"FF93", X"FFF8", X"FE6A", X"FF76", X"0228", X"0020", X"00A9", X"000C", X"00A1", X"00DD", X"005B", X"FF94", X"0079", X"FD5A", X"FEAF", X"009E", X"00A7", X"FF74", X"FFB5", X"FF8C", X"01E2", X"FB57", X"FF47", X"0486", X"00F4", X"0124", X"0385", X"001D", X"FFAB", X"012F", X"FFA9", X"00D0", X"0027", X"FF88", X"007B", X"FF65", X"FEF0", X"0029", X"0105", X"00C9", X"FF69", X"FAAC", X"FA24", X"F869", X"F92A", X"F9C9", X"FE68", X"FF2C", X"FFE8", X"00A2", X"01FD", X"0359", X"0201", X"FFA1", X"FDA9", X"FDC3", X"FC7D", X"FBD9", X"FD9A", X"FF4F", X"0053", X"00DF", X"0017", X"FFFE", X"003D", X"001D", X"0217", X"016C", X"0015", X"FF0F", X"FFF0", X"FE65", X"FE2A", X"FDEE", X"FF78", X"0221", X"0417", X"025B", X"02F7", X"035F", X"02D2", X"01E7", X"FE25", X"FC51", X"FC1F", X"FAC3", X"FC24", X"FF51", X"0080", X"0005", X"017C", X"0009", X"FECC", X"FDDC", X"FF11", X"FDE7", X"FF76", X"FFAB", X"FF11", X"FFDF", X"0045", X"0312", X"01DE", X"0405", X"057A", X"04D2", X"02BE", X"045B", X"0114", X"0058", X"FF8A", X"FE81", X"FFFF", X"FEC4", X"0193", X"0375", X"FFCC", X"FFC6", X"FFD2", X"0096", X"002C", X"FCDE", X"FEC0", X"FC2B", X"FE7D", X"FE45", X"FF30", X"FFD2", X"00A0", X"FFCB", X"0134", X"002E", X"003E", X"0263", X"00A4", X"0349", X"0217", X"0329", X"FFBA", X"014B", X"0378", X"02C9", X"0449", X"050D", X"FFDE", X"006D", X"FF0F", X"FC06", X"FE6F", X"FBC3", X"FC9D", X"FE4C", X"FDA8", X"FF7E", X"0049", X"00FF", X"FFB4", X"013B", X"0035", X"FFD6", X"00F8", X"FF99", X"FFC9", X"FE6A", X"000A", X"0089", X"FE4A", X"FF97", X"035C", X"0743", X"08FA", X"0692", X"026B", X"FFCC", X"038D", X"FA48", X"F994", X"FCB2", X"FE17", X"FCF0", X"FFA2", X"01B3", X"FF8C", X"FF4F", X"FF71", X"FEDB", X"00A0", X"0213", X"0190", X"0055", X"FF53", X"FFB1", X"00AB", X"01F1", X"002C", X"0125", X"026E", X"06C2", X"0897", X"04C1", X"02C9", X"009E", X"FDB7", X"F980", X"FBA9", X"FDA0", X"FF42", X"FF7D", X"0086", X"0156", X"00F2", X"FE11", X"009B", X"00AC", X"0088", X"02BA", X"034D", X"0058", X"FE2D", X"0019", X"0181", X"00EB", X"0189", X"01E0", X"020C", X"07A9", X"096E", X"04CB", X"021D", X"FEA9", X"FBA7", X"FE08", X"FBFA", X"FB77", X"FE2F", X"FF89", X"0216", X"0058", X"FF43", X"FD3A", X"001E", X"00CE", X"00BF", X"03E1", X"02C9", X"FEAE", X"FEE7", X"FE22", X"FEE6", X"0025", X"02D2", X"01C5", X"0327", X"0802", X"0D37", X"08F6", X"03AB", X"FDEB", X"FBED", X"F959", X"FB45", X"FDC5", X"FC74", X"FFC9", X"FF94", X"002C", X"FF67", X"FFEC", X"FFC7", X"0051", X"0336", X"07AE", X"0923", X"0188", X"FCFA", X"FD5B", X"FE21", X"FE51", X"FEBB", X"FDB3", X"027F", X"0A7F", X"0E25", X"09FD", X"037C", X"00B3", X"FBD6", X"FBB0", X"FCEF", X"00CC", X"FEE2", X"0077", X"FE2F", X"FEE6", X"FF9E", X"FF37", X"FEF7", X"01EB", X"0684", X"0975", X"0961", X"039A", X"FDB4", X"FFD5", X"FF9B", X"FCEF", X"FB00", X"F98B", X"FF1B", X"0706", X"0BCD", X"082B", X"020A", X"FDFC", X"FB54", X"F725", X"FC9F", X"FED0", X"000A", X"FEFE", X"FF6A", X"FF9D", X"0284", X"FFD1", X"FE5F", X"0224", X"06A5", X"0995", X"0798", X"012A", X"FD66", X"FEEE", X"FFDE", X"FF5C", X"FA49", X"F79D", X"F4FC", X"F590", X"FFD9", X"02AF", X"FDBA", X"007B", X"FDF7", X"FA0E", X"FC28", X"FD75", X"FD69", X"FE51", X"FF1F", X"FE4E", X"00E6", X"FDDD", X"FE74", X"0240", X"09D3", X"0831", X"05EE", X"0150", X"FD50", X"FF6D", X"FCE8", X"FE0A", X"F824", X"F4C0", X"F28E", X"F147", X"F6CA", X"FAE4", X"FDE2", X"01B2", X"FF99", X"FCFE", X"FC00", X"FC8E", X"FD72", X"FB4D", X"FC66", X"FDE8", X"FFFA", X"FE37", X"FFAF", X"0412", X"07A0", X"08FD", X"0466", X"FED3", X"FBB4", X"FC10", X"FAB8", X"F880", X"F9B3", X"F667", X"F503", X"F873", X"F980", X"FA31", X"FDFA", X"028E", X"028B", X"0453", X"FD2A", X"FB63", X"FBBB", X"FD29", X"FA5C", X"FBC1", X"FD0A", X"FC86", X"00CB", X"08D0", X"0A2D", X"0657", X"FE8D", X"FA17", X"F7E3", X"F93C", X"F921", X"F93C", X"F9A1", X"F95D", X"FB2F", X"FF0A", X"FB12", X"F95C", X"FCAB", X"FF06", X"03C0", X"054E", X"01A2", X"FF98", X"FE77", X"FD48", X"FA58", X"FCF9", X"FCEC", X"FDAF", X"0259", X"0922", X"072C", X"0142", X"F8D1", X"F722", X"F7B1", X"FA5A", X"F99D", X"F905", X"F8D2", X"FAAF", X"FF5A", X"027F", X"F8EB", X"F7C0", X"FEEA", X"FF12", X"02DA", X"00A5", X"02DE", X"03E0", X"001D", X"FF75", X"FDA8", X"FCDB", X"FBA7", X"FC2C", X"014F", X"0737", X"011E", X"FAA7", X"F5FD", X"F8E2", X"FA5C", X"FAA1", X"FCDF", X"FCA2", X"FD19", X"FE9D", X"0316", X"01CE", X"F80E", X"F6DE", X"FB2A", X"FDC6", X"FFFE", X"0313", X"0476", X"01FB", X"0029", X"0197", X"FE52", X"FE38", X"FFBF", X"FFB6", X"02A8", X"041C", X"FE63", X"FD7E", X"FCA2", X"FBE2", X"FBC8", X"FB22", X"FE06", X"FE73", X"FF02", X"00A0", X"03C9", X"0033", X"F966", X"F98B", X"FD71", X"0054", X"FA29", X"01CF", X"03D0", X"0149", X"01DB", X"FFD9", X"FEA3", X"FF8B", X"0209", X"0101", X"FED9", X"00CF", X"006B", X"FFE4", X"0094", X"FF74", X"FE6B", X"001C", X"00FB", X"00E3", X"0269", X"015C", X"034A", X"012E", X"F980", X"FA9B", X"0113", X"005F", X"FD38", X"FF8C", X"018E", X"01E3", X"005E", X"FFEE", X"0131", X"02F6", X"016B", X"01B6", X"FE55", X"FE9D", X"0203", X"0265", X"0279", X"01A6", X"043F", X"0422", X"03BD", X"04AD", X"033F", X"05B6", X"04F8", X"FDC7", X"FA34", X"FC04", X"FFD8", X"FFC6", X"FF56", X"FFB0", X"01AC", X"01E8", X"0016", X"0230", X"01B9", X"00D5", X"FF6E", X"FFC7", X"FFE6", X"00CA", X"027D", X"022F", X"0422", X"0462", X"057D", X"059A", X"03F4", X"064D", X"02F5", X"03B9", X"0089", X"FC85", X"F98F", X"FC1B", X"0078", X"0016", X"0076", X"0117", X"0205", X"02C5", X"FF51", X"00C0", X"010D", X"FDBB", X"FE23", X"FDA9", X"FF71", X"002D", X"014B", X"0337", X"011C", X"0414", X"046D", X"05BE", X"0449", X"060B", X"04C1", X"03C0", X"00B6", X"F95B", X"F9EF", X"00BB", X"0057", X"FE85", X"FE9A", X"0576", X"0792", X"05DA", X"01E4", X"0023", X"FEA8", X"FE88", X"FEAE", X"00DC", X"FF97", X"FFFA", X"0150", X"00A4", X"01FB", X"03EF", X"058A", X"0392", X"04B2", X"0474", X"0082", X"00EA", X"FF39", X"FD8C", X"FB89", X"0228", X"0133", X"0077", X"00D3", X"0202", X"0538", X"0369", X"FF8C", X"00A9", X"007F", X"01E9", X"0110", X"02D8", X"01C1", X"0281", X"0223", X"0389", X"0326", X"01DA", X"0289", X"04E8", X"03DB", X"0253", X"FD17", X"00A6", X"01C6", X"FE02", X"FD33", X"FCE8", X"0007", X"FF5B", X"0059", X"0186", X"FE57", X"FE9A", X"FD4B", X"FEE8", X"FDC9", X"0277", X"01B3", X"033D", X"0235", X"0308", X"02E3", X"008B", X"0016", X"0241", X"0430", X"0310", X"009E", X"FF37", X"FE90", X"0532", X"060E", X"05AA", X"FCE6", X"FD31", X"01E3", X"0084", X"0032", X"FFD9", X"FF71", X"FD1A", X"FC43", X"FA6D", X"FD36", X"FDB3", X"FEB0", X"FF70", X"0322", X"0062", X"FEFB", X"FEF5", X"FE05", X"FF85", X"FDB7", X"FCC7", X"FB98", X"FECB", X"00FD", X"FF74", X"00E3", X"FF99", X"007E", X"FFDC", X"0039", X"FFED", X"FFD6", X"FFAD", X"FF7E", X"FEFA", X"FDAC", X"FEAC", X"FDD3", X"FBBD", X"FF69", X"FF85", X"FF3B", X"FD1E", X"FB77", X"FBC6", X"FD69", X"F990", X"F6FD", X"FB0F", X"F940", X"FB13", X"FC0A", X"FD50", X"FEDF", X"FFDE", X"FFD3", X"FF55", X"FFCF"),
        (X"FE94", X"006F", X"0000", X"003E", X"00BD", X"FF84", X"FEAC", X"FFD5", X"FFEA", X"002B", X"FF31", X"FFCF", X"00BA", X"FFE9", X"FFA2", X"FF4B", X"FFE8", X"FF98", X"0018", X"00BF", X"0153", X"00B9", X"000E", X"00CE", X"006F", X"FFDF", X"0096", X"FFE0", X"0116", X"001C", X"FEAD", X"FF4A", X"FF96", X"00FD", X"0124", X"0207", X"FFFB", X"02E8", X"03B3", X"03CF", X"04D9", X"04CA", X"0275", X"0270", X"0508", X"03B3", X"0138", X"0281", X"0400", X"03F1", X"0345", X"0286", X"FE72", X"0295", X"FFA1", X"FF63", X"017E", X"0032", X"FF51", X"0172", X"0171", X"FEEF", X"0110", X"0362", X"0325", X"05EF", X"090E", X"0751", X"0947", X"0962", X"0978", X"07DB", X"080D", X"06B2", X"0881", X"076E", X"06A3", X"0475", X"05FB", X"0435", X"01EF", X"00B4", X"FFBA", X"FFE9", X"0119", X"004F", X"FDA4", X"FF9D", X"0070", X"02C4", X"02A3", X"0441", X"05D2", X"0754", X"0761", X"0913", X"0BD7", X"0B90", X"0E02", X"0CF9", X"0B80", X"09C9", X"0A18", X"0715", X"06C8", X"05C4", X"044E", X"05BB", X"05EF", X"037B", X"0279", X"002B", X"0159", X"FF18", X"FE96", X"006D", X"0036", X"02FB", X"0069", X"029B", X"0371", X"02C2", X"02C1", X"0396", X"048E", X"0500", X"07C3", X"0572", X"03A7", X"0583", X"059C", X"000B", X"FF2E", X"FFFA", X"FE44", X"0055", X"04B3", X"0869", X"0600", X"02F1", X"FEC6", X"00A5", X"FF82", X"FE4A", X"014C", X"FEC7", X"FEC8", X"005C", X"0182", X"FFB6", X"0007", X"0103", X"FF2B", X"0223", X"016B", X"0195", X"0232", X"0483", X"05BD", X"0475", X"0302", X"01B2", X"FE33", X"FE02", X"FFB9", X"070A", X"052E", X"02DF", X"009C", X"009F", X"00E6", X"FDBD", X"0037", X"FFC8", X"01B1", X"00CF", X"018E", X"FFFE", X"FFC2", X"FD96", X"FFE9", X"FFFC", X"001B", X"02B4", X"024E", X"0196", X"00EC", X"0333", X"0235", X"0088", X"FE85", X"FFDF", X"FF5A", X"0553", X"0169", X"03AD", X"0000", X"0120", X"0061", X"FCB0", X"001A", X"0159", X"027D", X"0382", X"01ED", X"0120", X"FFCF", X"FEC5", X"FF70", X"FECF", X"021B", X"0227", X"0189", X"00F0", X"0172", X"008C", X"00A4", X"FF74", X"FF34", X"FDED", X"026F", X"04A9", X"0002", X"044E", X"01E2", X"0285", X"0075", X"FE1F", X"FF81", X"FF5C", X"035F", X"011B", X"019E", X"024A", X"01BD", X"009F", X"0137", X"0100", X"0188", X"01B5", X"0263", X"0093", X"0216", X"0208", X"03BB", X"01FE", X"00B8", X"0235", X"05D4", X"04D7", X"0307", X"01B2", X"FF60", X"0293", X"0143", X"0022", X"008D", X"0164", X"01D9", X"0317", X"02EB", X"02EA", X"0328", X"01A3", X"012A", X"0060", X"0084", X"FE62", X"FE44", X"0060", X"0081", X"01FC", X"031A", X"041E", X"0264", X"056F", X"085C", X"0A6B", X"07AF", X"FF09", X"00A7", X"00A3", X"02E5", X"025C", X"01E6", X"0278", X"050A", X"04D2", X"0228", X"03F9", X"0314", X"0025", X"0010", X"0285", X"FEA6", X"F912", X"FBB3", X"FD41", X"0129", X"02AA", X"0273", X"02F0", X"03AC", X"0C61", X"09D4", X"07CF", X"0552", X"FFEE", X"FFDD", X"01AF", X"0354", X"FF52", X"010D", X"03A3", X"0362", X"02E2", X"FEEA", X"FFE3", X"FDFF", X"FD63", X"FE6D", X"00BC", X"FA55", X"F849", X"F863", X"FC89", X"FE4F", X"FF0F", X"FF51", X"0258", X"062B", X"0AFA", X"0CB3", X"0900", X"05B1", X"FDAC", X"FFA1", X"FD84", X"01CD", X"FFC6", X"FF59", X"02F5", X"028C", X"FE53", X"FD4B", X"FDD3", X"FC55", X"FD7D", X"FD65", X"FD9D", X"F8D7", X"F9C8", X"F978", X"F96A", X"FBEC", X"FDAF", X"FF7C", X"0172", X"04C3", X"06D3", X"0919", X"0772", X"05AA", X"008A", X"FE39", X"FD26", X"0197", X"FFF1", X"FCEB", X"FFD4", X"0132", X"FCB3", X"FD18", X"FA88", X"FE3A", X"009F", X"FE90", X"FBA6", X"FA3F", X"F9BB", X"FA68", X"FAD6", X"FC26", X"FD5E", X"FFA0", X"00A3", X"04E6", X"075E", X"0785", X"069C", X"051E", X"020F", X"0162", X"FFE3", X"0106", X"FE77", X"FB7E", X"FF6A", X"00FA", X"FDDE", X"FE5B", X"FD30", X"FFAC", X"0110", X"FE82", X"F9E8", X"FB00", X"FBBD", X"F9F8", X"F984", X"F935", X"FE76", X"022B", X"02D7", X"0402", X"05F4", X"08DB", X"053F", X"0384", X"0224", X"0139", X"FFFE", X"FFB6", X"017F", X"FE95", X"024A", X"0452", X"001E", X"001D", X"FFF7", X"0080", X"FF7B", X"FE0B", X"FB25", X"FC7F", X"FC8B", X"F9A6", X"FA45", X"FB5C", X"0251", X"049E", X"0302", X"030C", X"05BE", X"08DD", X"0865", X"0415", X"FF5D", X"FFAF", X"00B9", X"01C4", X"03E6", X"02C0", X"0560", X"0642", X"025A", X"0081", X"0080", X"0198", X"00FB", X"FDBC", X"FC7D", X"FBCB", X"FE14", X"FA7C", X"FEC1", X"023A", X"04B2", X"04FC", X"03B4", X"0642", X"075F", X"0959", X"092A", X"078C", X"02AF", X"0079", X"FE58", X"01D7", X"0447", X"06A3", X"0943", X"0B3E", X"0893", X"0397", X"038E", X"01DE", X"02BF", X"FF86", X"FBE0", X"FBBB", X"FE3B", X"0084", X"04BB", X"0633", X"0726", X"0731", X"0590", X"0805", X"0774", X"0805", X"07D1", X"041C", X"02F2", X"0017", X"FEA8", X"01A9", X"022A", X"0647", X"09E3", X"0C38", X"0918", X"08DD", X"0634", X"068B", X"0505", X"0306", X"005A", X"FEF9", X"03FD", X"0725", X"0857", X"0968", X"0909", X"0766", X"08A0", X"091D", X"0973", X"08A6", X"07A6", X"FF64", X"FE76", X"0033", X"0128", X"012E", X"020E", X"046D", X"0689", X"076F", X"0611", X"0655", X"07C0", X"0772", X"0672", X"04DB", X"027E", X"0287", X"052E", X"05A6", X"086B", X"08E1", X"08D1", X"0992", X"06D9", X"0A02", X"0A14", X"07D4", X"0410", X"0088", X"FD0B", X"00CD", X"0141", X"0342", X"068A", X"046D", X"04CF", X"02AD", X"02C4", X"0326", X"05DD", X"034C", X"0407", X"03C6", X"0527", X"0387", X"04E4", X"0339", X"034D", X"05EB", X"03DC", X"080A", X"06B7", X"0697", X"07F4", X"04DF", X"01F1", X"FFE8", X"0081", X"013B", X"FFAD", X"04DD", X"055F", X"0180", X"FDB4", X"FE17", X"0176", X"0035", X"00F9", X"0041", X"0215", X"0430", X"06AB", X"046F", X"02EC", X"01EF", X"01B6", X"032F", X"03CF", X"05A1", X"059D", X"060E", X"057A", X"0249", X"00B9", X"01F8", X"00FD", X"FF88", X"FF80", X"03A2", X"00D6", X"FEC8", X"FAAB", X"FC12", X"FF09", X"0025", X"FE22", X"FEFA", X"0263", X"0381", X"045F", X"0390", X"018D", X"0146", X"FF03", X"FE76", X"0018", X"00BE", X"03EE", X"04F9", X"021F", X"00F2", X"FF11", X"FDF4", X"003C", X"FF10", X"00E4", X"03D7", X"0426", X"006D", X"F9C1", X"FD8F", X"FD15", X"FE16", X"FF70", X"FE57", X"0099", X"0042", X"00D4", X"0246", X"015D", X"FD2A", X"FA4A", X"FE09", X"FCC6", X"0017", X"0020", X"FFFB", X"0113", X"FF0B", X"FEF7", X"FC39", X"00E8", X"0055", X"FF76", X"0260", X"0331", X"01D1", X"FAC9", X"FD35", X"FEFC", X"018C", X"0239", X"03C5", X"037C", X"04A5", X"0511", X"057D", X"0490", X"036F", X"0137", X"FED6", X"FE25", X"FEE8", X"FEB8", X"FEDF", X"FD96", X"013A", X"FF8E", X"FF5B", X"FFCD", X"00C7", X"FF97", X"0074", X"FBCA", X"FCCB", X"F9B4", X"FDB2", X"FE09", X"00DE", X"021E", X"00FF", X"0508", X"04E4", X"03C2", X"03F1", X"0454", X"0338", X"02E4", X"032D", X"0189", X"FFC7", X"FF70", X"FFA3", X"FD86", X"0092", X"0049", X"FF26", X"FEDC", X"016E", X"0030", X"0010", X"FEDA", X"FC21", X"F9E4", X"F9B4", X"FEF9", X"00D3", X"00D7", X"0203", X"02AB", X"01BC", X"033E", X"0081", X"028A", X"02CF", X"003B", X"0151", X"0082", X"00C4", X"0032", X"FFF0", X"FFB4", X"004C", X"007E", X"00C1", X"0058", X"FE57", X"0098", X"0192", X"000C", X"005B", X"01CF", X"01C8", X"02AE", X"03A7", X"026B", X"04C2", X"017F", X"0111", X"0602", X"03C3", X"02A3", X"05AE", X"0631", X"025C", X"FFF4", X"FF07", X"00FD", X"FF5B", X"FF65", X"FEA7", X"FF2B", X"FE96", X"FF4D"),
        (X"0135", X"000F", X"0092", X"FEBE", X"0056", X"0042", X"002B", X"FD48", X"FF93", X"FE5F", X"FF01", X"FFF5", X"0077", X"FFBF", X"0090", X"0035", X"01BD", X"008A", X"0049", X"0033", X"FF74", X"FFA1", X"FF13", X"0001", X"FF59", X"003E", X"FF1F", X"00F7", X"FFAA", X"0042", X"FEF4", X"00A5", X"002A", X"012E", X"021D", X"020C", X"047F", X"03BB", X"0279", X"04E6", X"041E", X"03E4", X"FC29", X"FDFA", X"01A9", X"033A", X"0329", X"03CC", X"02FE", X"024E", X"02B1", X"FFDC", X"FF4D", X"014D", X"FFE5", X"FFE7", X"FFB1", X"FF9F", X"001D", X"042A", X"032D", X"0106", X"00B3", X"0260", X"022A", X"011F", X"0299", X"0542", X"02DB", X"FD27", X"F96F", X"FBC4", X"0158", X"04DA", X"0510", X"02A6", X"0416", X"0219", X"005F", X"FFDC", X"FC95", X"FC18", X"00E4", X"FF42", X"FFCC", X"FF4B", X"00BF", X"021C", X"0196", X"FCBE", X"0091", X"01D7", X"0498", X"01EC", X"025E", X"03CE", X"046A", X"0351", X"0032", X"0233", X"00BE", X"04C4", X"04DC", X"0675", X"08A0", X"04A3", X"0182", X"FFAD", X"0163", X"00EA", X"01B0", X"FDF0", X"FF9F", X"FF33", X"FD32", X"02FE", X"FEF6", X"FFBA", X"0145", X"0193", X"FFAF", X"0236", X"02FE", X"0469", X"02B2", X"00B5", X"00C6", X"01B4", X"FF51", X"FEB6", X"007D", X"0138", X"FEA2", X"FF88", X"0289", X"0356", X"01EF", X"0486", X"FEEE", X"FD1B", X"FE2B", X"002E", X"0045", X"01C9", X"FC94", X"0186", X"026A", X"0155", X"00DA", X"0184", X"022F", X"012B", X"0062", X"01A6", X"0014", X"00CE", X"01B4", X"00AC", X"0292", X"0222", X"012E", X"020A", X"00BB", X"00EF", X"02DF", X"01A8", X"0136", X"FEC3", X"0046", X"00F4", X"FFC9", X"017D", X"FF65", X"01BF", X"01E7", X"FF17", X"0252", X"01F7", X"FFFD", X"FFF9", X"001D", X"00A2", X"00B6", X"FFF1", X"0146", X"037A", X"03BD", X"0289", X"0379", X"0135", X"FFB5", X"0066", X"03F2", X"0234", X"0486", X"FFC2", X"FFFA", X"0173", X"FDF9", X"021B", X"0123", X"02AA", X"FFFA", X"FE58", X"009C", X"00C9", X"FFF1", X"0116", X"00F2", X"FF12", X"0089", X"FEC2", X"003E", X"0199", X"02E5", X"02D0", X"0200", X"001C", X"FE90", X"000B", X"0113", X"04FE", X"01F7", X"0381", X"0060", X"FF56", X"FE26", X"019B", X"FCE4", X"FCA5", X"FA91", X"FC07", X"0074", X"003E", X"FDB8", X"FF6D", X"0012", X"FE43", X"FEE6", X"FF1E", X"0257", X"017B", X"03B6", X"01AD", X"0348", X"017C", X"0154", X"028E", X"02AF", X"0296", X"01D0", X"015F", X"FEE8", X"FF02", X"FFF0", X"FEB5", X"FDF1", X"F9CB", X"FE64", X"FDD4", X"FE2E", X"FE0B", X"FD98", X"FD99", X"FC05", X"FD1D", X"FF40", X"FF56", X"FF15", X"FF32", X"0172", X"0132", X"02FC", X"03CA", X"0539", X"0547", X"09FC", X"08B1", X"0391", X"04C7", X"FF06", X"FF46", X"0138", X"026C", X"FD49", X"FB4D", X"FCD6", X"FD84", X"FE83", X"FCC7", X"FC5E", X"FC69", X"FDE1", X"0083", X"00D2", X"FFCF", X"FDF8", X"FF08", X"00A9", X"00F6", X"01C7", X"01B9", X"04A5", X"0676", X"0CE5", X"0D8E", X"096B", X"0035", X"FF21", X"FEDB", X"FFF0", X"FC76", X"FBCE", X"FB7F", X"FBD4", X"FBB1", X"FDB0", X"FBB9", X"FD02", X"FE26", X"FF4C", X"023F", X"00CF", X"FD25", X"FDC0", X"FDDF", X"FE95", X"FFC4", X"FD19", X"FDD4", X"FD1B", X"03D8", X"09C5", X"0B47", X"0596", X"01CE", X"FF42", X"FE3F", X"FE2A", X"FCFE", X"FB90", X"FD92", X"FF59", X"FE42", X"FD88", X"FFA9", X"0416", X"02D0", X"03B3", X"05DD", X"FF53", X"F9DC", X"F98E", X"FA67", X"FC13", X"FBDE", X"F8D9", X"F651", X"F5F7", X"F9E4", X"FC72", X"FE9F", X"0263", X"FF19", X"0061", X"0025", X"FF03", X"FCC4", X"FC38", X"FF7C", X"FF86", X"0018", X"0164", X"0291", X"064D", X"0528", X"054F", X"018A", X"FCCD", X"F811", X"F806", X"F98B", X"FB3D", X"FA31", X"FA5E", X"FA72", X"FB46", X"FA92", X"FDD4", X"F7BD", X"FF99", X"FDBB", X"0285", X"00C2", X"0007", X"FD1C", X"FEE2", X"FFAA", X"002F", X"04B4", X"0562", X"060F", X"0729", X"041D", X"011F", X"FD28", X"FB75", X"FB2D", X"F76E", X"FA1B", X"FBE3", X"FD93", X"0212", X"031D", X"FF06", X"01BD", X"043E", X"FA52", X"F8A4", X"FEFD", X"00AD", X"0218", X"0005", X"FD11", X"0299", X"0197", X"028D", X"04EA", X"0621", X"05D2", X"0303", X"FD5E", X"FC9C", X"FDCE", X"F9D8", X"F9CF", X"FA43", X"FA1D", X"FE41", X"00BC", X"0643", X"0874", X"02DF", X"01A8", X"0639", X"FA4C", X"F986", X"FBFE", X"FE06", X"0030", X"0427", X"0245", X"0481", X"0784", X"0502", X"0290", X"0263", X"FB22", X"F974", X"F8AC", X"FC66", X"FAC4", X"F978", X"F99E", X"FBB9", X"FD81", X"00AF", X"02C3", X"06CE", X"0571", X"0527", X"0490", X"0327", X"FA49", X"F833", X"FE87", X"0131", X"0198", X"01D5", X"03DD", X"0520", X"0ABF", X"07DC", X"02FA", X"FBFD", X"F619", X"F670", X"F89C", X"F7DE", X"F7BB", X"F782", X"F9F9", X"FDD6", X"03DE", X"0368", X"056A", X"0461", X"0343", X"04C5", X"032B", X"010E", X"F832", X"F939", X"03EF", X"0052", X"FFF5", X"0264", X"053A", X"09C2", X"0B27", X"08B7", X"0415", X"FEA4", X"F85C", X"F964", X"F8AB", X"FB6B", X"FC51", X"FBF3", X"FE4F", X"0252", X"0587", X"03DE", X"0397", X"02BB", X"0324", X"0405", X"02ED", X"FF91", X"F784", X"FAD2", X"FBDF", X"0059", X"053A", X"04B1", X"061D", X"087C", X"08D2", X"06DB", X"02E6", X"056E", X"00CA", X"0014", X"00D6", X"01D3", X"000A", X"FF29", X"02B2", X"0329", X"02F1", X"02FE", X"02AC", X"00BF", X"040F", X"038A", X"01F5", X"FFDB", X"F683", X"FCAD", X"FE19", X"FF90", X"044B", X"05B3", X"060A", X"082F", X"071E", X"054B", X"0215", X"05A4", X"05EB", X"045A", X"0385", X"0390", X"02E2", X"0355", X"01ED", X"0216", X"0107", X"FF85", X"FEB3", X"FFCD", X"01E0", X"0333", X"04E9", X"FFB2", X"F8F5", X"FCCC", X"00A8", X"FFE5", X"0072", X"0449", X"0831", X"05F1", X"032A", X"0194", X"0165", X"02A1", X"FF75", X"01CD", X"0305", X"032E", X"0305", X"00EA", X"00FE", X"FF71", X"0016", X"FD84", X"FEDA", X"00AB", X"008E", X"0348", X"0279", X"FD5D", X"FCE2", X"0146", X"008E", X"0000", X"00E4", X"032C", X"0638", X"03E5", X"0009", X"001F", X"FF5E", X"00FF", X"012E", X"01BE", X"0333", X"02D8", X"00BC", X"00E2", X"013B", X"0013", X"002C", X"FE6B", X"00C6", X"FF4E", X"FEEB", X"00DF", X"02F0", X"FEBA", X"FE63", X"0338", X"013C", X"00A6", X"FF6D", X"0455", X"0854", X"0741", X"0624", X"0171", X"0158", X"00B8", X"037C", X"03B6", X"03C4", X"0179", X"0182", X"0044", X"0152", X"021C", X"FE20", X"FE99", X"FDCB", X"FF15", X"FDB0", X"FFEB", X"00F6", X"0175", X"FFF4", X"045D", X"0069", X"0037", X"008C", X"021B", X"06B9", X"082C", X"06CD", X"03AD", X"01BD", X"0022", X"006D", X"00C5", X"0234", X"01B1", X"0203", X"03CA", X"0220", X"0165", X"0349", X"0210", X"FDF6", X"FD9C", X"FE8A", X"FFF6", X"FFB3", X"017F", X"FD8E", X"FF38", X"00C5", X"FF69", X"FF91", X"01F1", X"0255", X"01FB", X"0191", X"FFBA", X"0058", X"FF5A", X"FFE4", X"0033", X"0218", X"021A", X"02DD", X"FF44", X"0105", X"0093", X"0330", X"01E4", X"0261", X"FF11", X"FE97", X"0334", X"0219", X"024E", X"014E", X"0013", X"0005", X"FF4C", X"0042", X"FFBB", X"FFBD", X"FE43", X"FD86", X"FA99", X"F8AE", X"F90D", X"F90B", X"FCA8", X"017B", X"02DD", X"FF89", X"FDF7", X"FE6C", X"FF75", X"0045", X"FF2E", X"020B", X"0205", X"013F", X"0055", X"FF89", X"00C3", X"00EC", X"007D", X"FEB2", X"FF48", X"00BE", X"FF58", X"FFB6", X"007F", X"FFF9", X"00C5", X"FE74", X"FE1E", X"FDD3", X"FF89", X"FF27", X"00FD", X"FD5D", X"F900", X"FAD7", X"FC63", X"FB46", X"FAFC", X"FA79", X"FD37", X"FE28", X"FD40", X"FD1E", X"0006", X"FEE2", X"000C", X"0013"),
        (X"0179", X"FFB1", X"00AD", X"FF1F", X"FF6D", X"FEF9", X"FFBE", X"0079", X"FF30", X"FE4B", X"FFCF", X"FFAA", X"0119", X"02B1", X"FFC0", X"FE98", X"0000", X"0076", X"FFC5", X"009F", X"015A", X"FF21", X"019E", X"FF87", X"0127", X"006B", X"010A", X"FFEF", X"00ED", X"0085", X"017C", X"004B", X"00B1", X"0116", X"0222", X"03F4", X"02CB", X"02CE", X"0242", X"0351", X"03CC", X"024B", X"024A", X"0201", X"0333", X"01B6", X"00B1", X"0261", X"0222", X"00BA", X"01F8", X"00B7", X"FFFF", X"FF4C", X"FFB3", X"006E", X"FF5E", X"FEFE", X"009A", X"00D2", X"FFF1", X"00C3", X"03F9", X"0635", X"0661", X"07ED", X"06F6", X"07E1", X"09BE", X"0A3E", X"0A54", X"068F", X"079D", X"03ED", X"022D", X"0203", X"010C", X"042B", X"0280", X"0406", X"01B2", X"0077", X"FF9C", X"FFC9", X"FFF4", X"FF9E", X"00D0", X"009E", X"FFDA", X"FF33", X"03D8", X"080A", X"087D", X"0952", X"095B", X"09ED", X"0BBA", X"0CB7", X"0AEB", X"07E7", X"0760", X"07BA", X"032C", X"01EB", X"0367", X"03DC", X"0353", X"01DC", X"015C", X"02EC", X"0074", X"0062", X"FE2C", X"FF6B", X"FF21", X"0078", X"FC96", X"FB8F", X"FEFC", X"FE4D", X"0100", X"0327", X"04CE", X"03C8", X"03E0", X"02BE", X"02CF", X"03A7", X"060B", X"04FA", X"00DC", X"0114", X"0387", X"00F0", X"FE6B", X"FB6F", X"FB9A", X"FB98", X"018A", X"039E", X"FF97", X"FF91", X"FFF3", X"FEB7", X"FB62", X"FB63", X"FBC0", X"FE34", X"00FF", X"01BF", X"004B", X"00D3", X"001F", X"FF90", X"0013", X"0175", X"03AA", X"02D8", X"025A", X"023D", X"FF97", X"0292", X"FE2D", X"FCB0", X"FDDD", X"FCE0", X"021D", X"0140", X"0071", X"0074", X"FECD", X"FE1A", X"F9BA", X"FE05", X"FE38", X"02A9", X"011C", X"0013", X"00DD", X"FFFC", X"FF9F", X"FE33", X"FE0C", X"01BE", X"FFF2", X"01BF", X"FF55", X"0054", X"FF06", X"011A", X"FEC3", X"FD2D", X"FC0C", X"FDE6", X"FD2E", X"0029", X"00BB", X"FDF5", X"FF13", X"FF1B", X"FE35", X"006B", X"013B", X"01A5", X"0033", X"FFEA", X"00A8", X"0151", X"0070", X"FEB9", X"FF9D", X"FFBD", X"0029", X"FFC8", X"00AD", X"FF95", X"FF6E", X"FFD1", X"00AA", X"0196", X"FD69", X"FE76", X"FE16", X"0062", X"FF53", X"03A8", X"FF8A", X"00CA", X"00CD", X"FFD3", X"015D", X"0020", X"FFF0", X"FEFA", X"0114", X"0256", X"0338", X"0081", X"00AD", X"008D", X"0165", X"000D", X"0170", X"00FE", X"0196", X"FFFC", X"01C7", X"02ED", X"FF5F", X"FDA6", X"FE60", X"FFAE", X"00DC", X"01A1", X"0060", X"02D0", X"0101", X"024B", X"FEF7", X"FEA0", X"FFE4", X"FEED", X"01D2", X"00B6", X"0173", X"FF4A", X"0136", X"011F", X"0111", X"01F7", X"023C", X"0094", X"0034", X"0058", X"0307", X"0200", X"FF91", X"FBD0", X"FE83", X"0193", X"00B9", X"033D", X"03AE", X"01DA", X"03D2", X"02B1", X"0210", X"019F", X"FF7C", X"01BC", X"0079", X"0194", X"012D", X"036B", X"04B4", X"04CD", X"0414", X"0187", X"01D1", X"0331", X"007F", X"00CC", X"00B3", X"00D4", X"FDB2", X"F8C6", X"FDCB", X"0314", X"003F", X"048B", X"0761", X"056F", X"04A9", X"0292", X"FF19", X"00A5", X"0074", X"02B2", X"02F3", X"0184", X"0493", X"0723", X"061F", X"025A", X"0217", X"00C2", X"011A", X"018B", X"FF55", X"00F3", X"FEA3", X"FEC1", X"FF94", X"FA8D", X"FD9D", X"025F", X"019D", X"03C8", X"085C", X"06CD", X"02B7", X"018F", X"FEA9", X"0081", X"007D", X"FEC1", X"FD79", X"FD14", X"FB23", X"F7D9", X"FB49", X"FDD0", X"0025", X"00C7", X"FF8D", X"FEE8", X"FEDF", X"FE06", X"FAD7", X"FDDB", X"0258", X"03D2", X"03BC", X"058E", X"FFDB", X"028B", X"066C", X"06F9", X"FD5E", X"FC94", X"FC4A", X"FCCB", X"FBFD", X"FDE4", X"FC54", X"F9CC", X"F7E4", X"F689", X"FA5E", X"FCF7", X"FEE2", X"FE03", X"FEAE", X"FEF6", X"FCD3", X"FD3F", X"FED0", X"FFF8", X"076A", X"0A4F", X"06C1", X"0311", X"0114", X"015B", X"047A", X"0467", X"FF73", X"FCCF", X"FA03", X"FB0A", X"FA64", X"FA40", X"FCE2", X"FDFC", X"FA2F", X"FDC7", X"FBB9", X"FCC4", X"FB3D", X"FDBC", X"0061", X"012B", X"FFE8", X"FF11", X"02CB", X"0358", X"0527", X"0744", X"0843", X"00D4", X"0149", X"FE9C", X"0209", X"03B1", X"0081", X"0014", X"FD95", X"FC06", X"FAEB", X"FCED", X"FC52", X"F9D7", X"FB31", X"FC35", X"FC82", X"FCE7", X"FCCE", X"FEA5", X"01DB", X"01BC", X"03EC", X"00DB", X"0137", X"01E0", X"0304", X"0A08", X"0116", X"023C", X"FFA2", X"FFEA", X"01C2", X"049C", X"05C3", X"0392", X"03E5", X"0202", X"FCE8", X"FBE6", X"FA2A", X"F7C4", X"F846", X"FC80", X"FBD3", X"FC4D", X"FE76", X"0097", X"00E9", X"0252", X"0366", X"00F3", X"0013", X"014E", X"0274", X"09E6", X"06B7", X"024D", X"0089", X"FED5", X"FDA1", X"04BB", X"0A54", X"0911", X"09F5", X"08B4", X"04F2", X"0489", X"FE46", X"FB9E", X"FF18", X"FE6D", X"FE4A", X"FDCD", X"00E9", X"028C", X"01A5", X"01F0", X"0461", X"019F", X"0314", X"03B1", X"06D7", X"0B4A", X"063B", X"01AD", X"01AB", X"0021", X"FE8E", X"0322", X"0A63", X"0B4C", X"0E64", X"0FD6", X"1076", X"0FA3", X"0CA5", X"09F3", X"0853", X"0591", X"049D", X"0111", X"018F", X"02CF", X"029D", X"02A5", X"01D0", X"0167", X"006E", X"0279", X"05EA", X"0A05", X"05A9", X"0129", X"010C", X"0446", X"00F2", X"01CD", X"0544", X"08AB", X"0D48", X"12FE", X"165D", X"1674", X"1488", X"1251", X"1197", X"0B35", X"065C", X"03D4", X"015F", X"0229", X"004E", X"0181", X"FED7", X"FD58", X"000E", X"0153", X"0258", X"04E1", X"01B6", X"FF63", X"FF51", X"01E6", X"FDFB", X"FB50", X"00AD", X"0360", X"062A", X"0B9E", X"0C8E", X"0D1C", X"0DAD", X"0CDB", X"0D4D", X"08A0", X"0650", X"017F", X"FF76", X"FF8E", X"010A", X"FF92", X"FD22", X"FC53", X"FE67", X"FD19", X"013A", X"FF4E", X"01A1", X"0157", X"FFBD", X"FEBD", X"FBB5", X"FE08", X"FA47", X"FD4A", X"FFED", X"0200", X"FEEE", X"01A4", X"FF65", X"0361", X"03FC", X"02AC", X"02B9", X"015F", X"FEE8", X"FE3C", X"FF5B", X"FE07", X"FCC7", X"FD02", X"FBFD", X"FCDF", X"FED5", X"FF34", X"013C", X"FF13", X"FFEC", X"00B8", X"FC7F", X"FC58", X"F964", X"FD27", X"FC28", X"FC84", X"FAAB", X"F921", X"F92E", X"FB14", X"FE4E", X"0023", X"FFF5", X"0121", X"0066", X"0011", X"0003", X"FF1F", X"FFA3", X"FE6C", X"FBCF", X"FA33", X"FE80", X"005D", X"0031", X"FFBE", X"FFD0", X"00A0", X"FAB4", X"F8D1", X"F806", X"F8D9", X"FB82", X"FAAE", X"F6F6", X"F9A9", X"F9FA", X"FA3C", X"FC83", X"FF3F", X"0072", X"00E9", X"01BC", X"00DA", X"026D", X"0192", X"FE92", X"FDA3", X"FA78", X"FA22", X"FD2B", X"FFD3", X"FEA9", X"004F", X"FF8B", X"FFF7", X"FF18", X"FB79", X"F943", X"FA0D", X"F9A5", X"F94C", X"FB4F", X"FA94", X"FA9B", X"FDCB", X"FEFD", X"0074", X"0034", X"020B", X"0301", X"FF35", X"0299", X"0277", X"001E", X"FC72", X"F898", X"F5D7", X"FE7A", X"01F4", X"02B4", X"FE7E", X"0096", X"FE64", X"FE58", X"012F", X"FFDD", X"FB1C", X"FAFE", X"FA6A", X"FD34", X"FC38", X"FC90", X"FF24", X"FD69", X"FDE6", X"0183", X"011A", X"0163", X"FF4D", X"021C", X"025B", X"FDCC", X"FBCB", X"FC01", X"F9A1", X"FC44", X"01C8", X"02C4", X"FF72", X"FEE6", X"0024", X"FEC5", X"FE87", X"F9A6", X"FC00", X"FC5C", X"FEA2", X"FF16", X"FE24", X"FEA0", X"FF23", X"009F", X"FE12", X"FF9B", X"0158", X"00F0", X"0236", X"0349", X"040E", X"FF17", X"0113", X"01C5", X"FE22", X"FEFD", X"FE57", X"FF6D", X"001F", X"FFEF", X"FF92", X"FFF6", X"FF68", X"FF02", X"FF0A", X"011A", X"FFDF", X"0312", X"FF89", X"FFAE", X"FE7C", X"FF42", X"047C", X"FF9B", X"FF95", X"01DD", X"02B0", X"00D2", X"0318", X"0147", X"0310", X"0388", X"025E", X"FF13", X"FE28", X"FF13", X"016F"),
        (X"FFF4", X"FF81", X"FF9A", X"001D", X"FFF9", X"0027", X"0097", X"FF2F", X"FFA8", X"FF49", X"00D6", X"FFD2", X"FF11", X"FC8C", X"014B", X"0044", X"FED4", X"FFA0", X"0021", X"00A0", X"008E", X"FFE1", X"FFA8", X"FF61", X"013A", X"0001", X"FF58", X"FF8D", X"FF53", X"0066", X"0016", X"0027", X"00A9", X"0008", X"FC30", X"FC5B", X"FB1B", X"FD20", X"FC8A", X"FD6C", X"FF36", X"FE67", X"FE53", X"0102", X"0417", X"FFBE", X"FC93", X"F996", X"F7A3", X"FC52", X"FCCF", X"FE22", X"FFDA", X"FE8C", X"0037", X"0038", X"FF72", X"00B1", X"FEFA", X"0191", X"FF28", X"FE13", X"FB53", X"F902", X"FB61", X"FC80", X"FAB4", X"F942", X"F926", X"FA5F", X"FAC6", X"FBD2", X"FCB3", X"FE61", X"FCB5", X"F937", X"FBBA", X"FA52", X"FA02", X"FC07", X"FDB7", X"FEEE", X"0140", X"FF8E", X"FF8A", X"001B", X"FEFB", X"FFB9", X"01EE", X"FF38", X"FC29", X"FA7B", X"FCFF", X"FC20", X"FC73", X"FD9D", X"FE24", X"FEF2", X"FE27", X"FD92", X"FCDC", X"FED9", X"FDDD", X"F867", X"F985", X"FAF0", X"FCB0", X"FD8B", X"FFEF", X"0255", X"0095", X"019C", X"FE6E", X"FF27", X"0089", X"FF03", X"FDA3", X"00C8", X"003E", X"FF5C", X"FE99", X"FF76", X"FF3A", X"02AD", X"0486", X"01AB", X"01A3", X"00FC", X"FFBA", X"FD8B", X"FC4F", X"FAE6", X"FBF3", X"FF0A", X"020E", X"00CD", X"035E", X"0472", X"02E3", X"00DC", X"FF38", X"FED9", X"FD72", X"01AB", X"0182", X"002B", X"FFFC", X"0057", X"FF8A", X"020B", X"0249", X"0589", X"0385", X"0282", X"03DA", X"02B4", X"0322", X"0039", X"FF18", X"FD79", X"0339", X"0855", X"09B2", X"0711", X"049A", X"04DD", X"02FA", X"FFAA", X"FFA4", X"FF63", X"0153", X"FF4A", X"008D", X"01C1", X"007C", X"0274", X"004C", X"0038", X"006B", X"FF59", X"0150", X"042C", X"01D1", X"00D4", X"FEEB", X"FE3F", X"FF40", X"01B0", X"0557", X"085F", X"0820", X"071E", X"061F", X"031A", X"036E", X"00EC", X"00B6", X"FE2B", X"FFCF", X"FE04", X"00A2", X"0391", X"02D7", X"00B7", X"017A", X"FD01", X"FDEE", X"FE08", X"0014", X"FF4A", X"00AA", X"FEF3", X"009A", X"FCCF", X"FFD7", X"03DB", X"03C2", X"048E", X"054D", X"02BF", X"05A3", X"0750", X"0174", X"0340", X"00E4", X"FCBC", X"FF50", X"FD65", X"000F", X"041D", X"0321", X"0096", X"FEAA", X"FE76", X"00B5", X"01F1", X"FFD1", X"FFE9", X"FF43", X"FF32", X"028F", X"02C4", X"043D", X"0525", X"065E", X"0398", X"0144", X"00D1", X"0369", X"03FF", X"033D", X"010D", X"FEED", X"FCDC", X"FDAF", X"FECA", X"FF9E", X"0382", X"01F0", X"0161", X"0028", X"0243", X"0505", X"01BB", X"0090", X"FF22", X"FFF0", X"FF55", X"031B", X"0541", X"05A8", X"0522", X"0357", X"0085", X"FF56", X"01E3", X"05E7", X"0941", X"058D", X"FE77", X"FFEB", X"FBCB", X"FD4C", X"00D4", X"FFB2", X"03D5", X"0198", X"00D8", X"00C1", X"03C3", X"0378", X"01E7", X"FFF1", X"FEC7", X"009C", X"02E7", X"046B", X"058A", X"0763", X"0311", X"007F", X"FD01", X"FD1C", X"023E", X"0939", X"0870", X"073C", X"FFF8", X"FFBD", X"FBC8", X"F6B3", X"FECD", X"FF00", X"02FC", X"01E2", X"00B7", X"FF08", X"0109", X"0161", X"FF66", X"FB56", X"FC89", X"000D", X"015A", X"009A", X"03BB", X"0287", X"00D2", X"FD4A", X"FB22", X"F976", X"FE4C", X"073D", X"0C3C", X"0806", X"0006", X"FDBE", X"FBA0", X"F710", X"FAE8", X"FECB", X"001C", X"FF39", X"FD24", X"FFA9", X"01C2", X"FF31", X"FDBE", X"FDA8", X"FDCF", X"00BE", X"FF8B", X"FF37", X"FFD1", X"02C2", X"017B", X"FB6F", X"F5CD", X"F649", X"F8BA", X"FFDC", X"068E", X"051D", X"01DF", X"00CA", X"FCF7", X"FA4E", X"FBE3", X"FE14", X"FE94", X"FB28", X"FC2F", X"FEF7", X"0185", X"FFD7", X"00EA", X"0235", X"03AB", X"004A", X"FA67", X"FD8A", X"01B7", X"0311", X"FE09", X"FAB8", X"F6E4", X"F7F9", X"FA0D", X"00AE", X"0820", X"0776", X"04A7", X"0207", X"FD94", X"FB54", X"FC11", X"FE13", X"FF4D", X"FBA4", X"FCE9", X"0000", X"FFA4", X"0010", X"0031", X"0511", X"02FD", X"00D8", X"FB5B", X"FE01", X"0174", X"00BA", X"FE30", X"FC81", X"FD1A", X"FE16", X"FDA9", X"0059", X"030D", X"0629", X"0279", X"005A", X"0057", X"FB0D", X"FF37", X"040D", X"01D7", X"FCAD", X"FDBF", X"0031", X"02E2", X"0105", X"00DF", X"04B0", X"0275", X"FCDD", X"FC91", X"FE64", X"0149", X"00FA", X"001A", X"FDEF", X"FE78", X"0052", X"013D", X"029B", X"03D9", X"05E9", X"00D2", X"FEDC", X"0079", X"014A", X"0082", X"040A", X"02F8", X"012D", X"FE4E", X"FF6F", X"021D", X"016F", X"01CD", X"02F2", X"FF29", X"FB1F", X"FC76", X"FF11", X"03D2", X"02A4", X"019A", X"0219", X"0135", X"02C8", X"0586", X"051F", X"046C", X"07FC", X"0275", X"FF79", X"FE7E", X"0278", X"030B", X"036C", X"0588", X"049A", X"0425", X"03D4", X"025C", X"FF8B", X"FFDD", X"0269", X"FDF3", X"F911", X"FBDE", X"FF63", X"04DC", X"0243", X"0346", X"019A", X"026F", X"0614", X"079D", X"067A", X"02FF", X"03B6", X"02AF", X"FCAE", X"FE2B", X"0190", X"03BB", X"0301", X"0848", X"0997", X"06BD", X"066A", X"0399", X"01A2", X"001D", X"FE79", X"FC02", X"F94E", X"FE13", X"0120", X"0058", X"00C4", X"FFE7", X"01D7", X"03A7", X"0705", X"06C5", X"0796", X"0236", X"FF7A", X"FF8B", X"FF87", X"FC44", X"FF95", X"058F", X"04E2", X"0672", X"076B", X"07BF", X"0869", X"04BF", X"0193", X"FD42", X"FBD5", X"FD49", X"FC27", X"FDBA", X"FF41", X"0152", X"0044", X"FE3F", X"020D", X"0376", X"06BF", X"08E6", X"0423", X"02D7", X"02E0", X"FF15", X"001B", X"0160", X"03B2", X"07A6", X"0723", X"085F", X"0798", X"083F", X"08EE", X"0606", X"00AF", X"FD88", X"F99B", X"FCD2", X"FA45", X"FD0A", X"FDC6", X"FE1E", X"00EB", X"02CF", X"0327", X"05F2", X"0739", X"095D", X"07CA", X"04AE", X"0267", X"FF00", X"FF8F", X"FF4E", X"027C", X"0277", X"03F6", X"06D6", X"05C8", X"0541", X"025B", X"0255", X"FEAD", X"FD35", X"FC7B", X"FAFD", X"FB19", X"FD6D", X"FDE4", X"FF0A", X"01CE", X"0253", X"0325", X"019F", X"0771", X"09E0", X"040B", X"0287", X"0130", X"FEE5", X"00C6", X"FF93", X"0275", X"0693", X"03D2", X"0527", X"05AF", X"0486", X"02D4", X"008D", X"0008", X"003A", X"0076", X"006A", X"017D", X"004F", X"0067", X"02F9", X"02B2", X"0376", X"0277", X"059B", X"07CB", X"0835", X"0342", X"026B", X"FE42", X"00A3", X"FFCC", X"00F7", X"0213", X"072F", X"0468", X"051B", X"056B", X"05DA", X"0505", X"0207", X"FFB6", X"02C0", X"01F1", X"02C2", X"027D", X"014C", X"017C", X"02B3", X"06AC", X"0713", X"07F1", X"0844", X"0817", X"07DD", X"03A9", X"0279", X"FE53", X"FEC4", X"020B", X"00CF", X"FE99", X"FFCD", X"FE9D", X"FD78", X"FF31", X"FF10", X"017A", X"FE03", X"FC14", X"FC22", X"FDA1", X"FF16", X"0075", X"0051", X"0419", X"04D3", X"0608", X"0727", X"07C2", X"0700", X"03DE", X"039F", X"04AD", X"FFF0", X"FFE7", X"0026", X"001F", X"00D7", X"015E", X"FF51", X"FF25", X"FD6B", X"FD7E", X"FD11", X"FD3A", X"FC40", X"FCF6", X"FBAA", X"FA57", X"FD34", X"FD16", X"FEB4", X"00EF", X"0199", X"035C", X"0262", X"0422", X"01B8", X"0030", X"0016", X"FD6D", X"006F", X"006E", X"0014", X"FFDB", X"003D", X"FF68", X"00E5", X"0124", X"0031", X"FBD9", X"FD79", X"FB5F", X"FCE8", X"FE0B", X"FD75", X"FFF7", X"FE7A", X"FB40", X"FC67", X"FD95", X"FCB0", X"FC55", X"FF07", X"0008", X"FFB0", X"FE23", X"FF7C", X"001F", X"FF49", X"00C7", X"FFFC", X"FF8F", X"FF45", X"000D", X"FEC4", X"FFB1", X"FE57", X"0056", X"0105", X"FFB2", X"FFC7", X"FF25", X"004D", X"FE2A", X"F831", X"FC5E", X"FDF2", X"FBC7", X"FB18", X"FCD3", X"FD7D", X"FE2E", X"FD7E", X"FB8C", X"FF2F", X"FF52", X"FF4B", X"0147", X"FE91"),
        (X"009A", X"0003", X"FFC8", X"FFEB", X"00E8", X"0030", X"00A8", X"0053", X"006A", X"FF3C", X"FFD1", X"00A1", X"00AC", X"00E7", X"0140", X"FED8", X"FFB9", X"0040", X"FF9C", X"FE96", X"022F", X"FE06", X"FEE2", X"0099", X"0136", X"0077", X"FF5E", X"FF38", X"0023", X"FF63", X"00C9", X"FF68", X"FF7E", X"FFF5", X"FFE8", X"FFE9", X"012E", X"0188", X"00C8", X"FEC6", X"FE8C", X"FF78", X"FEC5", X"FC07", X"FE54", X"0000", X"006F", X"00A8", X"FFA5", X"FFC5", X"00C3", X"FEFE", X"00AF", X"00FF", X"FF5B", X"0082", X"0088", X"003A", X"FFFD", X"FDF0", X"FF5A", X"00FC", X"0054", X"FF3C", X"02F2", X"0791", X"0617", X"055D", X"0480", X"0062", X"00E8", X"007D", X"FECB", X"FEE7", X"FF71", X"000E", X"01B9", X"00DB", X"001F", X"FE20", X"0376", X"010C", X"FF84", X"FF65", X"FFC2", X"003E", X"FCBC", X"FE1B", X"026B", X"0392", X"0677", X"0529", X"029C", X"0426", X"0473", X"02B3", X"0087", X"004A", X"FE8C", X"FD51", X"FECA", X"FEB9", X"FF4C", X"01BF", X"0198", X"00AE", X"0195", X"0103", X"0163", X"FFC0", X"01FE", X"FEF0", X"FF8E", X"FF61", X"FCD5", X"FC5E", X"0197", X"0356", X"0579", X"0374", X"05C2", X"04B6", X"056F", X"0335", X"02C5", X"FF60", X"FEDB", X"FBF6", X"FF9F", X"FF68", X"0015", X"0200", X"01E0", X"0161", X"018C", X"0379", X"005E", X"FFC0", X"FD10", X"0191", X"004B", X"0016", X"0182", X"FDE7", X"02C1", X"0011", X"02A1", X"0193", X"02E6", X"01B1", X"FF47", X"FBD3", X"FC1C", X"FBE6", X"FB57", X"FC46", X"FB67", X"FCA0", X"FDF4", X"FE47", X"FD68", X"FB94", X"FC56", X"017D", X"FF10", X"FD1E", X"0016", X"0321", X"FFB5", X"FF0B", X"FF0B", X"FC3A", X"0177", X"0040", X"FDB7", X"FE56", X"FBCD", X"FB90", X"F987", X"FB2E", X"FA51", X"FB19", X"FD49", X"FBD5", X"FE1C", X"FF72", X"FDB5", X"FD05", X"FC88", X"FB08", X"FBE8", X"FEAD", X"FDA0", X"FFDA", X"0111", X"01B5", X"FF9A", X"FD8A", X"0096", X"FABC", X"FD16", X"FB42", X"FA54", X"F92B", X"F8BF", X"F9DC", X"F92D", X"FABC", X"FB3D", X"FC74", X"FDED", X"FD4A", X"FC94", X"FE1D", X"FC52", X"FD80", X"FDB7", X"FDE4", X"FC59", X"FC1B", X"FCFC", X"FE9F", X"0193", X"00FC", X"FDDC", X"FE3E", X"FFC0", X"FBBD", X"FC1F", X"FB08", X"FA15", X"F843", X"F97D", X"FAD0", X"FA49", X"FD9D", X"FC5A", X"FD44", X"FEDA", X"FC91", X"FC08", X"FA1A", X"FD09", X"FD53", X"FD57", X"FE25", X"FB9F", X"FC12", X"FAF9", X"0051", X"FBBB", X"FB74", X"FD82", X"FD6B", X"FD28", X"FB29", X"FB17", X"FC57", X"FAE8", X"FA9A", X"FA19", X"FD3D", X"FEB4", X"FD5B", X"FE6E", X"FF58", X"FFCD", X"FD2E", X"FB2C", X"FB4F", X"FD99", X"FDE0", X"FFA9", X"FE66", X"FCF3", X"F892", X"F8E8", X"F889", X"F8AB", X"FD31", X"FEC2", X"FB7B", X"FB96", X"FA02", X"FC80", X"FE3E", X"FEA9", X"FE6A", X"FEEC", X"FFFC", X"FDC0", X"FEC0", X"FF56", X"FABD", X"F967", X"FA26", X"FB04", X"FC24", X"FC7F", X"FE4E", X"FC4F", X"FDE1", X"FC82", X"FA25", X"F712", X"F93B", X"F733", X"FBEE", X"0002", X"FCF5", X"F85F", X"FAC2", X"FD20", X"01CE", X"FF5B", X"FE3A", X"0027", X"FFAC", X"FE5E", X"FD2C", X"FBB6", X"F5E8", X"F619", X"F93A", X"FD2D", X"FDC4", X"FFA9", X"FF7F", X"FFA7", X"FF75", X"FC29", X"F9CC", X"F4EB", X"F800", X"F81B", X"FF5C", X"FF72", X"FD8C", X"FB0F", X"FB62", X"FF23", X"FDE7", X"FFDF", X"0072", X"01BA", X"00EA", X"024A", X"00DA", X"FFDB", X"FE5B", X"0048", X"02AE", X"002A", X"00CF", X"0241", X"02F4", X"0124", X"001D", X"FCF0", X"F975", X"F9AE", X"FC6E", X"FBD1", X"FD13", X"00AC", X"FD05", X"FA74", X"FDC4", X"0360", X"0137", X"033B", X"038C", X"02E1", X"02CC", X"054D", X"0625", X"05C9", X"05AB", X"067D", X"0409", X"02FC", X"0213", X"031E", X"02DF", X"019C", X"0164", X"FE6A", X"FE22", X"FC88", X"FEE4", X"FD86", X"01D0", X"FCF3", X"FE4E", X"FBBC", X"FF9A", X"0240", X"01A9", X"032F", X"0459", X"0583", X"0430", X"0424", X"078D", X"0640", X"0728", X"0516", X"0406", X"058D", X"03C4", X"01EA", X"020B", X"0143", X"FFD1", X"FE14", X"FF06", X"FC47", X"0134", X"035F", X"019D", X"FEE9", X"0094", X"FE2C", X"01B7", X"02A0", X"0189", X"0588", X"0435", X"0364", X"0242", X"03E0", X"0492", X"02EF", X"012D", X"0356", X"053F", X"057A", X"0476", X"02A9", X"01B9", X"FF6B", X"FFB1", X"FF8B", X"FDD0", X"FD93", X"021B", X"06AE", X"026E", X"FF4C", X"FECA", X"FB3B", X"FFD6", X"FFDD", X"0198", X"0495", X"0490", X"032C", X"0220", X"01D0", X"0390", X"FFCE", X"015E", X"05C7", X"050B", X"069F", X"0575", X"0322", X"0080", X"00EF", X"021D", X"FF72", X"FF05", X"FF42", X"04F6", X"0624", X"02E7", X"0070", X"FED0", X"FE43", X"FC90", X"FCF8", X"0070", X"0335", X"063C", X"0607", X"01CD", X"051B", X"014B", X"FF3D", X"02F5", X"055A", X"075B", X"053D", X"023A", X"024F", X"0070", X"FF52", X"012D", X"003B", X"0024", X"FF0B", X"0598", X"041E", X"0172", X"FF1D", X"FEF7", X"FDDA", X"FF0E", X"0076", X"FF1F", X"FFBB", X"0584", X"04E3", X"049D", X"02A5", X"01D4", X"02D3", X"0531", X"0695", X"06D2", X"053B", X"01E4", X"035E", X"016C", X"FFA9", X"0051", X"FF36", X"0256", X"048F", X"0641", X"01E8", X"0415", X"00A2", X"FD88", X"FA7B", X"007C", X"00C8", X"FF74", X"FEF8", X"FFF7", X"0104", X"FFCD", X"01B3", X"031F", X"00BD", X"0233", X"0382", X"03D9", X"0446", X"02B2", X"01B1", X"00A8", X"00AE", X"0044", X"FF38", X"034F", X"04C9", X"0716", X"0500", X"0284", X"00D8", X"FE71", X"FD8B", X"01D6", X"0312", X"FDA8", X"FC05", X"FCBC", X"FD0B", X"FC8D", X"FC95", X"01C5", X"009C", X"012A", X"010B", X"01AE", X"0254", X"0091", X"00FC", X"012D", X"006B", X"FECA", X"00B0", X"0179", X"068C", X"0A32", X"024F", X"FE16", X"FF70", X"035D", X"FF97", X"013B", X"000D", X"FD73", X"F812", X"F9DE", X"FB25", X"FB06", X"FB95", X"FB32", X"FBB3", X"FEA8", X"FD49", X"FCB8", X"FD44", X"FD9D", X"FD90", X"FCF4", X"FD3E", X"FE24", X"FF84", X"02F1", X"0817", X"09D9", X"02B0", X"0019", X"007C", X"01BC", X"0103", X"0399", X"027B", X"FC73", X"F932", X"F90B", X"F901", X"FAFF", X"FADD", X"F9EC", X"FBA7", X"FAF1", X"F952", X"FA05", X"F9E1", X"F948", X"F9D4", X"FB9E", X"FB44", X"FF58", X"FEC8", X"0400", X"06A8", X"0637", X"FFE2", X"FF78", X"00A7", X"FFFE", X"0126", X"FFE3", X"FE33", X"FF39", X"FAB3", X"FBF2", X"FBA1", X"FB97", X"FB31", X"F9F8", X"F91E", X"FAA8", X"F98F", X"F89F", X"F6FB", X"F924", X"FAE3", X"00ED", X"FFED", X"01D0", X"00F3", X"01EF", X"066B", X"04FE", X"03D9", X"FFCD", X"FFEA", X"FF80", X"FEDE", X"FBF8", X"FE9A", X"FE7D", X"FEFF", X"0082", X"FF4F", X"FDB8", X"FC9D", X"FB79", X"FB84", X"F973", X"FB85", X"FAA1", X"FCDE", X"FDB0", X"015E", X"0191", X"0329", X"057C", X"02AD", X"03CC", X"0159", X"039A", X"01BD", X"FFDE", X"FEB7", X"FF67", X"025E", X"FCC1", X"FF7F", X"0374", X"0664", X"0467", X"038E", X"0245", X"0134", X"00FA", X"FF8A", X"FF25", X"0103", X"FFED", X"01C5", X"0181", X"021C", X"03E7", X"09FD", X"07A5", X"024A", X"025E", X"FF36", X"0005", X"FF4B", X"FEE6", X"FF22", X"FF38", X"010A", X"00C2", X"0578", X"0574", X"063F", X"051B", X"014A", X"0086", X"0271", X"00A2", X"01B0", X"011A", X"0290", X"0065", X"FFE1", X"0018", X"002F", X"0055", X"0545", X"0375", X"007A", X"02AA", X"0079", X"FF82", X"0009", X"FF27", X"00DE", X"00F3", X"018D", X"FFF2", X"FED5", X"FDCE", X"FFE6", X"FEA2", X"FC92", X"FC2A", X"FC4B", X"FEE3", X"004D", X"FAF4", X"0039", X"014D", X"FCA4", X"FD01", X"FF1D", X"FFD9", X"00FB", X"FE70", X"FE83", X"FC9F", X"FFE8", X"007D", X"FECF", X"0066"),
        (X"FFF2", X"FFC6", X"FEFD", X"FFAA", X"FE0C", X"FFCF", X"004A", X"FFEB", X"FF79", X"0035", X"00B5", X"00C5", X"FEDF", X"FEBC", X"FC94", X"FF14", X"0147", X"0026", X"FF48", X"FF83", X"FEAE", X"FEF9", X"017C", X"FF74", X"000C", X"FFE0", X"0037", X"FEEB", X"FFCE", X"0102", X"FFB5", X"FFC5", X"FFDB", X"FF76", X"FC72", X"FDF0", X"FD33", X"FD02", X"FD4B", X"FB5C", X"FB13", X"FBDA", X"0018", X"FAA1", X"F96E", X"FBDC", X"FB9C", X"FB65", X"FA74", X"FEC6", X"FE40", X"FE75", X"00C0", X"0006", X"00C5", X"FFDF", X"FFDB", X"FF46", X"FFD4", X"FEA2", X"FC3A", X"FE9C", X"FC15", X"F91C", X"F7F0", X"F4A9", X"F5F3", X"F617", X"F712", X"F768", X"F89C", X"F55E", X"F6A5", X"F6CC", X"F862", X"FBA4", X"FB9A", X"FACC", X"FA57", X"F9DD", X"FC37", X"FC9E", X"FF35", X"00DA", X"0031", X"0065", X"FD36", X"FCA9", X"FD8B", X"FF5F", X"FCFD", X"FD30", X"FC9F", X"FA74", X"FDAF", X"FBF9", X"FA99", X"FA15", X"FB8E", X"FBB2", X"FA4F", X"FC4E", X"FEB5", X"FD99", X"FFB3", X"FE70", X"FE9B", X"FFA9", X"FA68", X"FC4D", X"FD36", X"001B", X"FFE1", X"00E1", X"FE6E", X"0010", X"0161", X"02D9", X"FFE4", X"0202", X"0217", X"014C", X"031C", X"027B", X"FF75", X"FEAF", X"00CF", X"FFD4", X"00D3", X"FE86", X"FFC4", X"0029", X"FD7F", X"FD09", X"FDAF", X"FD7D", X"02EC", X"010A", X"02A6", X"FE6E", X"FF35", X"FFC4", X"FFD6", X"FDEC", X"01DA", X"0088", X"FFDE", X"FEF5", X"FDFF", X"FF5F", X"FF5E", X"01F0", X"FF73", X"FE71", X"FF48", X"FF6F", X"FF62", X"007A", X"0031", X"029C", X"0268", X"FE6B", X"FF22", X"FE3D", X"024B", X"05BD", X"00D8", X"FF25", X"FFBF", X"0226", X"004A", X"FFED", X"025E", X"FE6D", X"FDE3", X"FBE0", X"FDD4", X"FD36", X"0037", X"FFD2", X"FFF0", X"FE6C", X"0130", X"02CF", X"0050", X"025D", X"02B5", X"01FA", X"017C", X"FE8A", X"FE3C", X"0182", X"0213", X"0737", X"0329", X"FF6D", X"FF33", X"0162", X"0004", X"002D", X"0249", X"FE17", X"FD76", X"FCE6", X"FE70", X"FE72", X"FF96", X"FEBC", X"FF2D", X"FFBA", X"FE80", X"0165", X"019B", X"000D", X"FE60", X"FE55", X"00C5", X"FD36", X"FCCB", X"FE27", X"005A", X"049F", X"0356", X"FED3", X"FE9D", X"F96E", X"FCF9", X"000C", X"FEBD", X"0004", X"FFEB", X"FF78", X"002C", X"FCE2", X"FECE", X"FEE7", X"FFC1", X"FD25", X"FBEA", X"FB6A", X"FDEE", X"FB69", X"FD80", X"FDEF", X"FE0D", X"FE41", X"FF6F", X"FC56", X"0403", X"09E4", X"089F", X"0395", X"FED3", X"FB37", X"FC88", X"FDB9", X"FED3", X"FEC6", X"00F5", X"FFBE", X"FD48", X"FECF", X"FD77", X"FD05", X"FC4C", X"FA60", X"F793", X"F6F4", X"F951", X"FA85", X"FAEF", X"FBEA", X"FEBC", X"00E6", X"0164", X"FFDE", X"0159", X"0796", X"06B3", X"003D", X"FE73", X"FA58", X"FA07", X"FF94", X"00E9", X"00B3", X"00E7", X"00E4", X"FEB1", X"FC83", X"FD0C", X"FD11", X"FDDE", X"F835", X"F4D5", X"F457", X"F73E", X"FAF5", X"FE20", X"FD6D", X"FFA3", X"FF03", X"0080", X"0239", X"0224", X"05CD", X"03C8", X"0278", X"FF6E", X"FB71", X"FC57", X"01BB", X"0443", X"047A", X"034E", X"FF41", X"01EA", X"01CD", X"0266", X"04FF", X"06AD", X"0432", X"FFEF", X"FDD7", X"FFD3", X"0074", X"00E2", X"0342", X"0207", X"FEE7", X"FF36", X"FF87", X"027F", X"0725", X"0790", X"009F", X"FF62", X"FB60", X"FC29", X"02B3", X"057B", X"053F", X"03D9", X"0223", X"03A0", X"042C", X"0695", X"08FA", X"0C9A", X"0E59", X"0A64", X"0744", X"05A1", X"0367", X"0225", X"02A7", X"01A2", X"0157", X"0049", X"00D1", X"FDE0", X"FE6A", X"FF83", X"FC2A", X"FF56", X"FE02", X"FB91", X"0491", X"07B6", X"04EC", X"0258", X"0381", X"04BA", X"0317", X"0361", X"0652", X"0956", X"0B8B", X"09BD", X"0848", X"0928", X"061D", X"063D", X"050E", X"01D3", X"00EE", X"FF8A", X"F9C9", X"F735", X"FAD8", X"FB48", X"FBAC", X"FFF0", X"0329", X"FC73", X"05C5", X"08E3", X"0457", X"049B", X"031D", X"0347", X"0063", X"FF88", X"0272", X"0447", X"05B3", X"05DB", X"059E", X"06E1", X"06A6", X"01D5", X"03B0", X"0003", X"FDE9", X"FA3E", X"FA7A", X"F89B", X"FA01", X"F81D", X"FB8F", X"0069", X"002F", X"FEBC", X"0762", X"064A", X"03BB", X"02E2", X"01E6", X"01C8", X"FFD1", X"FD4C", X"FE75", X"03ED", X"0288", X"0300", X"04EF", X"0400", X"0197", X"019D", X"024F", X"0098", X"FF11", X"FEA3", X"FB6C", X"F9DF", X"F73D", X"FBEB", X"FD24", X"FEB4", X"0343", X"01DC", X"0866", X"02DA", X"FEDA", X"0197", X"0129", X"005A", X"FF6B", X"FCF7", X"0044", X"048B", X"0176", X"00AD", X"0416", X"0231", X"0072", X"0109", X"01B7", X"00C9", X"FDEC", X"FF45", X"FFD9", X"FCD5", X"F3A1", X"F819", X"FC7F", X"FFE3", X"016B", X"02C6", X"07A4", X"0202", X"FDF7", X"FF3B", X"00B6", X"FE6B", X"FE8B", X"FECA", X"FF64", X"0271", X"0069", X"024B", X"0417", X"0258", X"0126", X"02D4", X"01BA", X"0145", X"0054", X"0217", X"FFDA", X"FB00", X"F0DE", X"F741", X"FB34", X"FE3C", X"0127", X"01C8", X"05C0", X"02AF", X"00E2", X"00E2", X"FDBD", X"FDA3", X"FD48", X"FECD", X"FE11", X"FE8E", X"FEAF", X"FE70", X"0179", X"02CE", X"01BB", X"016C", X"0444", X"02AE", X"020E", X"025C", X"FF3B", X"FA65", X"F180", X"F778", X"FC35", X"FE80", X"FB76", X"0221", X"06C4", X"02ED", X"0342", X"FFC4", X"FCCC", X"FC1C", X"FB9D", X"F938", X"FBAF", X"F9C3", X"FB7D", X"FBDB", X"0027", X"01C6", X"03CE", X"04BA", X"042F", X"0329", X"0255", X"02BB", X"FF85", X"F9A7", X"F373", X"F8F5", X"FC6A", X"FFFA", X"FE13", X"0314", X"0407", X"0314", X"008F", X"FFC7", X"FE48", X"FD31", X"FB19", X"FA5C", X"F95B", X"F8F9", X"FB85", X"FB8A", X"FF0F", X"0344", X"061E", X"0455", X"0306", X"0275", X"02D9", X"0213", X"FE2E", X"F939", X"F796", X"FC95", X"0026", X"FF9F", X"FFE0", X"033E", X"04C7", X"0359", X"FEC2", X"0070", X"FE9D", X"FDF9", X"FC5E", X"FC68", X"FC22", X"FABD", X"FAED", X"FBE5", X"FD9A", X"0034", X"01DB", X"037F", X"013A", X"0135", X"0011", X"0100", X"FC8C", X"F8F0", X"F941", X"FA2E", X"00A7", X"FE2D", X"FFBD", X"03A3", X"0584", X"060C", X"FAE6", X"FD5A", X"FBD0", X"FB9E", X"FB25", X"FDB4", X"FD92", X"FE6E", X"FE14", X"FD6E", X"FD8B", X"FF28", X"02E9", X"0260", X"0137", X"006C", X"0023", X"FFC6", X"FDDB", X"FB5E", X"FC32", X"FE74", X"FF4A", X"0146", X"FF61", X"0379", X"07D9", X"0394", X"FFB8", X"FBAC", X"FD0B", X"FE77", X"FEED", X"00D4", X"FEC4", X"FDA1", X"FF29", X"FDCB", X"FD1B", X"FF18", X"00F9", X"02EC", X"02A6", X"00BC", X"0308", X"0205", X"0347", X"FBB8", X"FE18", X"FE1E", X"00E4", X"00A6", X"0115", X"01B4", X"0823", X"0381", X"FFF0", X"01BA", X"0299", X"0265", X"00FF", X"01FE", X"0034", X"FFE6", X"FF03", X"FDCC", X"FCD2", X"FFEE", X"FDAD", X"FF1E", X"02F0", X"0276", X"0356", X"0487", X"0431", X"FBE3", X"FCDC", X"FEE6", X"0164", X"FF69", X"FF95", X"027B", X"FF8D", X"00FD", X"010A", X"021A", X"0380", X"01B1", X"01B0", X"034E", X"FF66", X"000A", X"00B5", X"FF0F", X"FDCC", X"FD93", X"FC0E", X"FF5B", X"01B0", X"0541", X"03B4", X"037C", X"053A", X"FF2D", X"FF8B", X"000B", X"015A", X"FED8", X"0097", X"FF5A", X"013B", X"048F", X"003F", X"02C0", X"0254", X"003C", X"FE0D", X"FD40", X"FE64", X"FEBF", X"FFC2", X"FBF7", X"F9E3", X"FB52", X"F7EB", X"F936", X"F904", X"FFA8", X"00C4", X"FD5C", X"005E", X"001F", X"FF3B", X"FFE7", X"00E8", X"0131", X"FEAE", X"00D2", X"006A", X"FEFA", X"FE11", X"FE50", X"0138", X"FDD8", X"FD1E", X"FEC0", X"FEBD", X"FDD4", X"F812", X"FE15", X"FCA3", X"F97D", X"F667", X"FB89", X"FC8F", X"FEDB", X"FC81", X"FF7C", X"FBDF", X"FF53", X"0148", X"FF1C", X"00EF"),
        (X"005E", X"FF1C", X"0004", X"0019", X"00B7", X"FEED", X"FF4F", X"001D", X"FEB0", X"FFA7", X"0047", X"000A", X"003C", X"FF1C", X"0108", X"0024", X"FF85", X"FFF2", X"01A7", X"FF93", X"FE2B", X"FFF9", X"0055", X"00F1", X"FFED", X"FF92", X"FFD2", X"0121", X"002D", X"0019", X"0072", X"00BB", X"FF01", X"FEF3", X"FE1D", X"FD46", X"FC26", X"FA9A", X"F9FF", X"F74A", X"F86C", X"F982", X"FEA5", X"FC1D", X"FA6D", X"F931", X"FC76", X"FBB4", X"FC1F", X"FB20", X"FB42", X"FF05", X"0038", X"016B", X"0042", X"FF45", X"FE86", X"01E2", X"FE83", X"FD61", X"FCAB", X"FF42", X"FB2A", X"F9C9", X"F973", X"F4AE", X"F465", X"F3E7", X"F30F", X"F43A", X"F5CC", X"F54D", X"F5D7", X"F7E3", X"F716", X"F967", X"FAA9", X"FAA9", X"FC50", X"FAB3", X"FD4A", X"FD7E", X"004F", X"FF75", X"FFE4", X"FF61", X"0232", X"FCB2", X"FD3B", X"FD74", X"F944", X"F67E", X"F4BF", X"F507", X"F376", X"F05B", X"EE95", X"EFD9", X"EFB2", X"F151", X"F491", X"F839", X"F998", X"F6C2", X"FA16", X"F8A4", X"FCB5", X"FEDA", X"FB69", X"FD17", X"FD9F", X"FE73", X"0034", X"FE89", X"02ED", X"FF20", X"FECB", X"FB66", X"FA5D", X"F9F9", X"FA98", X"FA55", X"FB1D", X"FA1C", X"FA34", X"FA57", X"F8E9", X"F9F7", X"FAAB", X"FBC2", X"FAE3", X"009D", X"00B8", X"00ED", X"01F6", X"0245", X"FBFA", X"F773", X"FD5E", X"FDF6", X"0095", X"FFB4", X"0226", X"0188", X"FDF7", X"01B8", X"039A", X"0198", X"FF12", X"FE77", X"0027", X"0140", X"00DC", X"FF1B", X"FFDE", X"FF19", X"FE5C", X"FB0C", X"FCC7", X"FCD5", X"FDED", X"FF75", X"0245", X"02DE", X"01E3", X"FBBB", X"F9F4", X"FDC6", X"00AC", X"FE12", X"FE21", X"016F", X"FD8C", X"FFAD", X"024F", X"016E", X"FF41", X"0087", X"015D", X"01A2", X"00FE", X"00C2", X"FFBC", X"FF58", X"FFFF", X"005E", X"FE47", X"FDCC", X"FEB5", X"0040", X"019A", X"FEDB", X"FE44", X"FCC9", X"FD35", X"FE00", X"0177", X"FE22", X"FF82", X"047C", X"FE13", X"FE8B", X"FEB4", X"FF0C", X"FEC4", X"FF4F", X"FFE3", X"0109", X"00D1", X"01B2", X"FF67", X"FEDB", X"01CF", X"00CC", X"FF90", X"00B8", X"0027", X"0017", X"FFD2", X"0008", X"FB07", X"FA5F", X"FF7D", X"FCFA", X"FE58", X"0199", X"0125", X"0181", X"FFBE", X"FE15", X"FEAA", X"FE95", X"FF80", X"FFBB", X"FEF2", X"FF9A", X"FDD2", X"002F", X"FDD1", X"0025", X"FE96", X"00D8", X"027A", X"FDBE", X"FFB6", X"FD27", X"FD94", X"FB50", X"F9E9", X"F9F2", X"FE40", X"FD6E", X"0073", X"014C", X"FF35", X"00AC", X"FD30", X"FDBE", X"0044", X"0146", X"0094", X"FF9A", X"010E", X"0120", X"00A2", X"FF3C", X"0090", X"019E", X"035D", X"048A", X"0337", X"FF3E", X"FEAF", X"FD3D", X"FB5D", X"F7C7", X"F6B5", X"F713", X"FB55", X"FFC6", X"FE93", X"0103", X"FF53", X"FE1C", X"FCED", X"FE6F", X"FFF9", X"01FB", X"00DD", X"012C", X"016C", X"02B9", X"FECA", X"FFF8", X"FF54", X"0435", X"056B", X"046A", X"0304", X"01CE", X"007E", X"FF91", X"FE23", X"F4ED", X"F392", X"F698", X"FA4D", X"00F5", X"FF60", X"0107", X"010B", X"FF2B", X"FE1F", X"01AB", X"00E7", X"03D4", X"0381", X"02E3", X"04E5", X"0403", X"FFF7", X"FD92", X"00F7", X"0495", X"0512", X"0597", X"0385", X"FFB0", X"02F4", X"0289", X"001B", X"F63D", X"F0ED", X"F285", X"F956", X"FFA0", X"0232", X"FFD9", X"017A", X"FE66", X"01DF", X"014C", X"0568", X"0515", X"04E3", X"0458", X"023C", X"00A6", X"FD1F", X"FD0F", X"0163", X"047F", X"0549", X"04BA", X"051A", X"03D9", X"051F", X"06E0", X"02A3", X"FB8E", X"F283", X"F5F0", X"F879", X"006C", X"0042", X"0178", X"02C4", X"0172", X"0571", X"03A4", X"057B", X"03D1", X"0479", X"00ED", X"FFE7", X"FC5B", X"FBE6", X"FD70", X"031F", X"03BA", X"046D", X"0444", X"045C", X"052B", X"065F", X"0736", X"002B", X"F8F1", X"F56C", X"F758", X"F7C2", X"FCE6", X"FD66", X"FFA8", X"0129", X"050A", X"06A8", X"02C3", X"03FB", X"0356", X"0334", X"FD63", X"FB26", X"FA46", X"FDD5", X"0116", X"0306", X"0413", X"023E", X"057D", X"056C", X"0595", X"0403", X"0007", X"FEED", X"FB0F", X"F61C", X"FA1A", X"F97A", X"FD90", X"FD83", X"FE6C", X"0031", X"056C", X"04DE", X"0158", X"00AF", X"01C6", X"008E", X"FBA7", X"FA62", X"FC09", X"FF67", X"020A", X"01D6", X"0107", X"037B", X"02DB", X"0348", X"018B", X"00CA", X"FE31", X"FD6A", X"FDA5", X"F6F7", X"F76F", X"FAF7", X"FE8C", X"00D5", X"FEB4", X"0029", X"00B0", X"001A", X"004B", X"FEEB", X"019D", X"FF31", X"FB42", X"FB6F", X"FDE2", X"007F", X"0300", X"042E", X"00BB", X"01DE", X"038C", X"008D", X"FF49", X"FEA3", X"FEB4", X"FE39", X"FA1C", X"F915", X"F547", X"F940", X"FD24", X"0007", X"0189", X"0083", X"FB1E", X"FDD7", X"FBA8", X"F902", X"FC8C", X"FD12", X"FCAC", X"FC0C", X"FD9F", X"0336", X"0629", X"044C", X"0261", X"FE72", X"FE29", X"FD2C", X"FC2F", X"FDA8", X"FBBA", X"FA2C", X"F72B", X"F83B", X"F650", X"FAD3", X"FB06", X"01F8", X"010B", X"0062", X"FBA4", X"FB00", X"F979", X"F679", X"F79B", X"FB54", X"FC72", X"FB37", X"FE67", X"02A4", X"0568", X"02E3", X"FF24", X"FA95", X"FB01", X"FA4C", X"FAFE", X"FA77", X"F84E", X"F626", X"F251", X"F3C5", X"F8D5", X"FF7B", X"016A", X"0176", X"FFDC", X"FEA3", X"FBCF", X"FA40", X"F6D2", X"F78D", X"F926", X"FB1B", X"F8B5", X"F9A4", X"FB87", X"FF7A", X"00D9", X"0094", X"FD61", X"FE05", X"FAFB", X"FA31", X"F97C", X"FB1E", X"F727", X"F40E", X"F301", X"F557", X"F9E3", X"FED1", X"0221", X"FF6D", X"FE86", X"FC5F", X"F7EC", X"FAB4", X"FB67", X"FB2A", X"FAA6", X"FB59", X"FAA4", X"FB6E", X"FBDF", X"FD6F", X"FE47", X"FF66", X"FCD5", X"FFE7", X"FDE4", X"FBCB", X"FAEA", X"F856", X"F8E1", X"F7EE", X"F690", X"FB9A", X"FE43", X"FD2D", X"FF14", X"0062", X"FF76", X"FA68", X"F7D6", X"FAC0", X"FF9E", X"00CE", X"FD84", X"FD9C", X"FDC9", X"FE1A", X"FBF5", X"FAF6", X"FC10", X"FDDA", X"006B", X"0221", X"FFBB", X"FE75", X"FCE3", X"FC6C", X"FBB3", X"F789", X"FAC7", X"FDE6", X"FDBE", X"FE1D", X"01C0", X"0087", X"FFF5", X"FB00", X"FA27", X"FD0C", X"04C7", X"02AD", X"FF5E", X"FF53", X"FE6E", X"FF4D", X"FCE6", X"FDA4", X"FD3F", X"01A7", X"022B", X"027A", X"028E", X"025A", X"0150", X"FE2C", X"FE06", X"FD15", X"FE43", X"FFBA", X"FFE2", X"0379", X"014E", X"009E", X"FFCA", X"FC71", X"F889", X"FDF6", X"02B6", X"01F9", X"00C2", X"FE1D", X"FC06", X"FE6C", X"FD7F", X"FDC1", X"FDE1", X"FFC2", X"0115", X"02C1", X"0347", X"030D", X"014A", X"01B5", X"028D", X"01C6", X"FEFC", X"FE85", X"00BB", X"0320", X"0052", X"FFE7", X"FF45", X"FDEC", X"FACC", X"FE3D", X"03AC", X"018E", X"FDC9", X"FB29", X"F96A", X"FC31", X"FA50", X"FA8E", X"FB1D", X"FC68", X"FD53", X"FC94", X"FF73", X"00A8", X"015C", X"0312", X"03CC", X"0297", X"0085", X"FE4C", X"FD35", X"FEA9", X"013E", X"FE53", X"0032", X"FEC4", X"0006", X"00D2", X"0377", X"0137", X"0078", X"00C0", X"FF63", X"FC1D", X"FD4A", X"FFDC", X"FC9B", X"FCF4", X"F9EF", X"F898", X"FA5D", X"FDCF", X"FEC7", X"01D3", X"036B", X"010C", X"FF2E", X"FF48", X"FE33", X"FEFE", X"00B6", X"009D", X"FEBE", X"FFD3", X"FF42", X"0021", X"0454", X"08F5", X"09D0", X"08C5", X"078C", X"0573", X"0327", X"00CD", X"01B0", X"02EA", X"01F9", X"FEC9", X"00BF", X"006C", X"FFEC", X"016A", X"FFDC", X"01BB", X"020B", X"0232", X"FE44", X"00C4", X"FEAE", X"FEFD", X"0073", X"003A", X"00B0", X"FF56", X"0030", X"00CB", X"00E3", X"003A", X"029F", X"004D", X"FF55", X"0000", X"01E7", X"04EB", X"043B", X"0244", X"0244", X"02FA", X"03C2", X"0261", X"04DA", X"0394", X"027C", X"0017", X"0135", X"0115", X"004D"),
        (X"FF36", X"0065", X"FFE3", X"FFDB", X"0003", X"FF35", X"FF04", X"004A", X"0150", X"0026", X"FF54", X"0057", X"FEEE", X"FECD", X"FF7E", X"FFE6", X"FFA3", X"00D4", X"005B", X"FF60", X"FF14", X"00F4", X"0195", X"0010", X"FF3B", X"FF3C", X"FF97", X"013E", X"FE35", X"0137", X"FFEA", X"FF64", X"FF68", X"FE9A", X"FD3D", X"FCDA", X"FCB5", X"FB86", X"FE06", X"FC99", X"FD87", X"FD09", X"002C", X"FCCC", X"FB43", X"FDE2", X"FC43", X"FAEF", X"FBF8", X"FD7C", X"FD93", X"FE6F", X"0037", X"006F", X"FF42", X"00BE", X"FEA3", X"009A", X"0027", X"FEC6", X"FF66", X"FE15", X"FA87", X"F9E7", X"F837", X"F6DE", X"F7FB", X"F9B3", X"F7E3", X"F935", X"F9D0", X"F978", X"FDFD", X"FCFC", X"FC90", X"FF2D", X"FECE", X"FEF8", X"FFEF", X"FB0A", X"FEEF", X"00C8", X"0000", X"FF66", X"006A", X"009E", X"FF49", X"FDC5", X"FE6D", X"0117", X"FF00", X"FCA8", X"FC2E", X"FBDA", X"FB2A", X"FF10", X"FDDB", X"FD28", X"FCC3", X"FCA5", X"FD18", X"FFBA", X"0086", X"0053", X"FD8F", X"FD3E", X"FC79", X"FC76", X"FCED", X"0217", X"005D", X"000E", X"0017", X"FFB6", X"0188", X"008A", X"00DF", X"00C1", X"FF10", X"FF19", X"FF7F", X"FF40", X"FE1D", X"00A9", X"00EE", X"FF43", X"FDCF", X"FF01", X"FF30", X"FFD9", X"FEBA", X"009D", X"FF04", X"FECB", X"FE2C", X"FCAD", X"FFC1", X"0387", X"04FC", X"FEB8", X"0113", X"0104", X"FCA5", X"0148", X"0093", X"015F", X"0226", X"027F", X"00DA", X"00F1", X"FFBD", X"017F", X"01E8", X"0096", X"003B", X"FF7B", X"00B8", X"00F6", X"FF29", X"FD5A", X"FDE0", X"FC57", X"FE6C", X"FDDB", X"FC8B", X"03CE", X"0225", X"FDA2", X"FF34", X"019B", X"0187", X"025A", X"0233", X"044A", X"045E", X"02BD", X"03EC", X"03DC", X"0223", X"02A7", X"01E7", X"03C1", X"03D1", X"052F", X"0408", X"0623", X"0338", X"02FA", X"030A", X"01B1", X"02D2", X"03E8", X"FFE0", X"00F4", X"016F", X"0134", X"FF12", X"0160", X"005F", X"05CF", X"045F", X"057D", X"0585", X"0390", X"0428", X"03B8", X"0112", X"FFAA", X"0261", X"0460", X"0465", X"0509", X"0765", X"065B", X"06F8", X"0546", X"0522", X"041D", X"0344", X"07E2", X"00E4", X"0018", X"0187", X"00BF", X"0256", X"FDF3", X"FE5B", X"0709", X"0527", X"0382", X"03EC", X"0502", X"054D", X"0278", X"FE7E", X"FF75", X"FFE0", X"03EB", X"02AD", X"03E2", X"0703", X"03C1", X"073F", X"0724", X"0371", X"04AB", X"040F", X"0107", X"01D0", X"FFB0", X"0409", X"011C", X"00C6", X"012C", X"0030", X"03F2", X"0545", X"01EF", X"02EF", X"06D1", X"01DB", X"0036", X"007D", X"FFCA", X"0256", X"0261", X"FF3B", X"FF45", X"020E", X"0302", X"0475", X"0633", X"021B", X"FF96", X"025E", X"028D", X"FFBD", X"FEDF", X"0072", X"FF8D", X"0036", X"00DF", X"02BB", X"0423", X"0340", X"00FD", X"0285", X"01FE", X"0111", X"03FD", X"019D", X"0277", X"037F", X"00E3", X"FE61", X"FF0A", X"0110", X"0286", X"05BD", X"04DD", X"018D", X"00E9", X"01FF", X"FF05", X"FA73", X"FA23", X"FDE1", X"0208", X"FFA7", X"011E", X"03BF", X"02BC", X"012D", X"00C6", X"02CC", X"0295", X"04AA", X"0368", X"0664", X"0610", X"04C8", X"03CF", X"0097", X"00F0", X"01FE", X"045D", X"03B9", X"03CF", X"0138", X"FDDF", X"00B7", X"FC1E", X"FB75", X"FA9E", X"03A1", X"FF98", X"FFB6", X"00CB", X"02B0", X"063A", X"02B3", X"036D", X"05A3", X"0771", X"0532", X"08EE", X"072B", X"0461", X"0464", X"03B8", X"FFFA", X"00DE", X"0293", X"026E", X"0428", X"04DF", X"01AC", X"FF88", X"FFD5", X"009F", X"0003", X"FF4B", X"03EF", X"FDC2", X"005C", X"0289", X"012C", X"FF6F", X"04A8", X"0759", X"072A", X"054A", X"0457", X"058B", X"0368", X"007B", X"00D1", X"FD68", X"FD39", X"FE23", X"031F", X"02E6", X"0463", X"0392", X"03A5", X"007A", X"FEED", X"FC9B", X"FF5F", X"00B9", X"FD83", X"FCE8", X"0093", X"031A", X"0022", X"FDD7", X"0540", X"0338", X"01A6", X"01C9", X"0069", X"00F1", X"FF59", X"FF68", X"FDB7", X"F9EB", X"F8F0", X"FD97", X"003A", X"04E1", X"046D", X"027D", X"01FD", X"0138", X"FF7E", X"FF23", X"FF5A", X"FB97", X"FB97", X"FDDC", X"FFCA", X"01A1", X"00F5", X"FC91", X"0127", X"0122", X"FF2B", X"0032", X"00D3", X"00B4", X"00A1", X"FDE6", X"FB4F", X"F8D0", X"FA56", X"FB5B", X"FE90", X"02F3", X"028A", X"01DC", X"00C3", X"0173", X"FFEC", X"0084", X"FCB6", X"F97F", X"FE91", X"FD6A", X"0108", X"02F1", X"FFA5", X"FCF9", X"FE0A", X"FC0B", X"FB27", X"FE2A", X"02C7", X"FE4A", X"FBB1", X"FAE8", X"FBBE", X"FA43", X"F7CA", X"FB87", X"FF25", X"0184", X"01F5", X"00C4", X"00F8", X"FF8C", X"01CF", X"FEF4", X"FEC5", X"F872", X"FA8D", X"FCC2", X"FE9E", X"00C5", X"FF35", X"FE9A", X"FFE7", X"FC12", X"FAC1", X"FE3F", X"FF57", X"FD62", X"FBDA", X"FC04", X"FC16", X"FA91", X"F787", X"FCD5", X"FF38", X"0249", X"012C", X"FFAF", X"FF8F", X"FE47", X"00ED", X"FFB1", X"FC3B", X"F8AF", X"FCD8", X"FCAB", X"0085", X"0087", X"007A", X"FEE2", X"FFE7", X"FE32", X"FC9A", X"FCB6", X"FCE7", X"FD02", X"FC64", X"FC00", X"FA64", X"FA87", X"F96F", X"FD3A", X"FFFC", X"FDB0", X"011F", X"FF11", X"0103", X"0059", X"FE7A", X"FBEC", X"F83F", X"F693", X"FD34", X"FB67", X"FFC3", X"0192", X"FED7", X"000D", X"FEF9", X"01DA", X"FED4", X"FCB6", X"FBB8", X"FA2E", X"FA6D", X"F958", X"FB28", X"FB20", X"FC8F", X"FD9F", X"FEED", X"FE56", X"FD83", X"FEEB", X"FCA6", X"FD4C", X"FDE0", X"FB59", X"FA7B", X"F41D", X"FAA3", X"FD36", X"0018", X"0279", X"017D", X"FFC7", X"FE07", X"02B7", X"FF84", X"FE0B", X"FAFB", X"FA5D", X"FB4E", X"F9AF", X"FB19", X"FD65", X"FCCA", X"0017", X"FEEE", X"FD70", X"FCD9", X"FC2A", X"FC79", X"FD59", X"FCF8", X"FC37", X"F78C", X"F971", X"FBAC", X"FF66", X"FE86", X"FF83", X"0077", X"FF56", X"FC74", X"0002", X"0031", X"FF74", X"FDB1", X"FB8D", X"F973", X"FBB6", X"FCE6", X"FE53", X"FEA6", X"017B", X"0005", X"FC8A", X"FB3D", X"FAEF", X"FD15", X"FD14", X"FF62", X"FB90", X"F8B0", X"F767", X"FD12", X"FFAF", X"FF7C", X"FFA6", X"0036", X"FCFF", X"FADE", X"FC75", X"002B", X"028E", X"01E1", X"00E0", X"0083", X"02FC", X"048C", X"055F", X"03B8", X"00E5", X"01C4", X"FFE4", X"FD9D", X"FC98", X"FC49", X"FF30", X"027A", X"FF09", X"FCAF", X"F9DB", X"FD77", X"004F", X"001D", X"FFA4", X"0033", X"0568", X"01F7", X"FDD1", X"0087", X"06E5", X"05C3", X"0488", X"08F4", X"0866", X"05DC", X"0892", X"07A9", X"06BD", X"04CC", X"05BD", X"0362", X"FF2A", X"0101", X"02B3", X"0067", X"01BB", X"0263", X"FD98", X"FD39", X"00E8", X"015D", X"0005", X"0209", X"051C", X"05AC", X"0365", X"048B", X"079C", X"059A", X"065C", X"0832", X"0929", X"0761", X"0A6C", X"0B42", X"098A", X"0ABA", X"05D7", X"04AD", X"0428", X"03D0", X"0291", X"0487", X"0562", X"FC20", X"FC41", X"FC48", X"FF89", X"FF9F", X"FF04", X"008A", X"01FB", X"04FB", X"060E", X"05CC", X"061A", X"07BB", X"0951", X"083A", X"09EB", X"079C", X"0A5B", X"0C2A", X"0B9C", X"0AF6", X"09AD", X"083C", X"08EB", X"058E", X"03B2", X"041C", X"02F8", X"0057", X"FE5A", X"FEEB", X"011D", X"005A", X"FFB3", X"0091", X"01CF", X"01A2", X"0287", X"0379", X"0463", X"047C", X"03EF", X"0481", X"0511", X"0560", X"0675", X"06A6", X"06F2", X"065C", X"04BB", X"05D3", X"054F", X"05AA", X"032C", X"032F", X"012F", X"0006", X"FEF1", X"FE62", X"FE7C", X"00CE", X"002C", X"FEF9", X"00D7", X"01C4", X"0033", X"00B4", X"00C5", X"FF77", X"FFFB", X"010D", X"0142", X"0247", X"0208", X"00EC", X"00B9", X"00A4", X"0181", X"0321", X"FFD5", X"007A", X"00BA", X"02C1", X"FEC8", X"0032", X"FF1D", X"FE4D", X"011B"),
        (X"0030", X"FEED", X"00E7", X"FF07", X"00F5", X"FE93", X"0031", X"006D", X"FF14", X"00DE", X"FFC2", X"0075", X"00FB", X"0089", X"FF37", X"FFF9", X"0045", X"011A", X"FFF2", X"000E", X"00BF", X"FFDA", X"0059", X"FF88", X"00DB", X"00A7", X"FE62", X"0002", X"0014", X"FEF1", X"01D6", X"FE98", X"FF91", X"0062", X"FE84", X"FF8D", X"007F", X"0196", X"011C", X"FFD0", X"FEFA", X"FEDE", X"0006", X"FDCF", X"FF0B", X"FF09", X"00C5", X"FF8B", X"0197", X"00FF", X"00F9", X"FEFF", X"000A", X"FF2C", X"00DF", X"0137", X"FFA0", X"FF20", X"00A4", X"FD9C", X"FFD4", X"01D3", X"030D", X"00EE", X"052E", X"0784", X"057C", X"02BD", X"FFB9", X"FEEB", X"012B", X"01A8", X"0370", X"056D", X"0618", X"0606", X"03A5", X"04E3", X"0467", X"032C", X"00BC", X"003C", X"0036", X"FF6B", X"004C", X"0136", X"FD5E", X"FF97", X"017D", X"FD99", X"FFD8", X"FFAA", X"FFA6", X"009C", X"FF93", X"FB6A", X"F91C", X"FA8B", X"F984", X"FD44", X"FF36", X"00FE", X"044A", X"0518", X"0480", X"06C7", X"0492", X"055D", X"00F5", X"0007", X"00CA", X"0057", X"0024", X"00FD", X"0043", X"FC6F", X"FCD6", X"FC3B", X"FCBD", X"FD8A", X"FDB4", X"FF1F", X"FE70", X"FCBF", X"FC71", X"FA9E", X"FF7F", X"FFC2", X"0225", X"0458", X"0594", X"0631", X"08AA", X"0A53", X"0733", X"036A", X"0279", X"016E", X"0239", X"01A1", X"00E5", X"000A", X"FDBA", X"FC8D", X"FB78", X"FA35", X"FB5A", X"FD75", X"0144", X"0183", X"0032", X"FF88", X"FE3D", X"0108", X"00F7", X"025B", X"01EA", X"0691", X"063B", X"05C6", X"08FC", X"0BDE", X"0A7D", X"092F", X"05BD", X"05CB", X"046F", X"01A5", X"FF58", X"FE91", X"FDB3", X"F9E2", X"FB36", X"FAF6", X"FB8E", X"FDC6", X"FEB0", X"01E8", X"FDDC", X"FEDA", X"FF1B", X"FD60", X"0009", X"FFF2", X"00A4", X"01CE", X"017F", X"05F2", X"060A", X"06BE", X"08F0", X"090F", X"09F8", X"0691", X"04A3", X"035B", X"FE25", X"FE4B", X"FE10", X"FA6B", X"F92E", X"FB13", X"FBF8", X"FD97", X"FDF0", X"FEB4", X"FDA9", X"FD11", X"FA7E", X"FCF7", X"FDB0", X"FEBC", X"FF93", X"FE91", X"005E", X"0069", X"031F", X"065E", X"054B", X"0705", X"0B7B", X"06F1", X"046C", X"0176", X"FFCB", X"FDFC", X"FAD5", X"F9B4", X"F7F7", X"FB2F", X"FCF3", X"FB9F", X"FF58", X"FF3C", X"FE5F", X"FF14", X"FC78", X"FD83", X"FAB2", X"FA0B", X"FD15", X"FC1D", X"FD33", X"0031", X"003B", X"0463", X"0161", X"04B7", X"080E", X"06C0", X"0755", X"03E7", X"FF5D", X"FDDA", X"F989", X"F95D", X"F934", X"FD5E", X"FEA1", X"FE46", X"0085", X"0155", X"0212", X"03FA", X"0205", X"FC61", X"F5F3", X"F5E1", X"F9BD", X"FA3F", X"FD00", X"FF65", X"FE9B", X"0098", X"FE16", X"01AE", X"0684", X"0795", X"073E", X"024C", X"FF53", X"FD6B", X"F842", X"F8C1", X"FBCD", X"FE6A", X"0072", X"00E3", X"0625", X"0618", X"068E", X"054E", X"0520", X"FCB9", X"F8E8", X"F9E1", X"F904", X"FB41", X"FCD5", X"FD9A", X"FB6A", X"FBC4", X"FB7E", X"023F", X"09AC", X"0909", X"07D7", X"FF99", X"FFEC", X"FB8A", X"F97D", X"F8EF", X"FC6E", X"0142", X"0243", X"0145", X"05ED", X"040B", X"0376", X"0177", X"020C", X"001A", X"FEF8", X"FF94", X"FE9E", X"FC7F", X"FC15", X"FB14", X"FA00", X"FB52", X"FBBE", X"0204", X"0A99", X"0B6C", X"057B", X"FEA1", X"FF8A", X"FF43", X"FA07", X"F939", X"FEC9", X"0117", X"000A", X"007C", X"0127", X"012C", X"003E", X"0117", X"03F3", X"0383", X"0144", X"0211", X"009B", X"00C4", X"FF7F", X"FF79", X"0001", X"FEFF", X"FE47", X"01E6", X"052D", X"0365", X"03F4", X"FD02", X"FF78", X"FFF2", X"FA95", X"FB80", X"FE34", X"FF2B", X"0208", X"0141", X"FFEE", X"00B4", X"FFE9", X"0339", X"04BF", X"035C", X"0104", X"0333", X"027B", X"02B3", X"016B", X"026D", X"00FA", X"FEAF", X"FE67", X"0177", X"016E", X"0229", X"02F0", X"0328", X"02B3", X"FEAB", X"FB16", X"FE28", X"0092", X"FFF4", X"00BB", X"0202", X"00F1", X"0047", X"02B5", X"0455", X"0498", X"03E6", X"0136", X"0146", X"01FC", X"0181", X"FE45", X"FEFC", X"0145", X"FC5E", X"FBC0", X"FECD", X"FF7D", X"02FA", X"03A6", X"03EC", X"017B", X"FE5F", X"FC22", X"0079", X"FF63", X"FED2", X"FFAD", X"006B", X"0256", X"0272", X"0328", X"03D3", X"0352", X"0371", X"026B", X"01A6", X"024E", X"FFA3", X"FDB7", X"FB58", X"FBD9", X"FCBA", X"FA09", X"FBC1", X"FF4B", X"0653", X"033D", X"0030", X"FE55", X"FD16", X"FC4F", X"FD71", X"FD2C", X"FF1A", X"016D", X"006C", X"02A3", X"FEBE", X"02E6", X"0336", X"03A3", X"04BB", X"028A", X"0469", X"0240", X"FF87", X"FD50", X"FCE5", X"FD58", X"FC31", X"FCAC", X"FCE3", X"0094", X"09C6", X"04C4", X"FFB6", X"FEC3", X"FE1C", X"FF48", X"FD4F", X"FE0D", X"0154", X"03D4", X"02F7", X"0307", X"02B2", X"020F", X"0545", X"06E9", X"04B6", X"0445", X"0265", X"017B", X"001D", X"FEA1", X"FC08", X"FE70", X"FC9E", X"FB58", X"FF57", X"0518", X"06F0", X"018D", X"FCA7", X"FCE0", X"FF0C", X"FDB7", X"FA80", X"001E", X"0299", X"04F4", X"0716", X"0475", X"04E3", X"034C", X"0814", X"08ED", X"083B", X"0395", X"009A", X"0063", X"FE89", X"0094", X"FEC4", X"FE61", X"FB5E", X"FC01", X"0293", X"0931", X"08A9", X"FFD3", X"FE88", X"004D", X"FBB8", X"FB9F", X"FD04", X"FFE8", X"0447", X"0562", X"03C8", X"0410", X"03CA", X"046F", X"073F", X"042D", X"0262", X"FF5C", X"01AA", X"00CE", X"FE66", X"FEFF", X"FECF", X"FE4D", X"FF07", X"01CE", X"0505", X"0686", X"0525", X"034A", X"FD51", X"FF1A", X"FE07", X"FD08", X"FBD4", X"002F", X"030D", X"03C7", X"046B", X"0437", X"01E6", X"02FE", X"02E5", X"0264", X"0087", X"FDB6", X"FF2C", X"FEFC", X"FF77", X"FFC5", X"FF3F", X"FEA7", X"02CB", X"02F6", X"064B", X"0715", X"027A", X"0045", X"FE67", X"FFFC", X"012E", X"FAC9", X"FDA8", X"0085", X"029B", X"01A8", X"02DF", X"053E", X"0558", X"02C1", X"01AE", X"FFB4", X"FFC9", X"00D3", X"FE0C", X"FE1F", X"FE5B", X"FEAB", X"0088", X"0106", X"03D7", X"06DB", X"080B", X"0833", X"02FA", X"01FD", X"FF7E", X"00C3", X"FFE4", X"FD6D", X"FD13", X"FF9E", X"FF93", X"00C8", X"0168", X"02DD", X"0351", X"FFC0", X"012F", X"FF9D", X"FF2D", X"FF52", X"FC0D", X"FE7B", X"FE95", X"FF9F", X"FF19", X"02BB", X"0641", X"07E7", X"08D3", X"082E", X"05B7", X"FF7D", X"FFEE", X"FEFC", X"003F", X"FD2F", X"FCD0", X"FC00", X"FD0E", X"FDC8", X"FDEE", X"0343", X"00C7", X"FDB6", X"FD70", X"FEB6", X"FD08", X"FE03", X"FE1D", X"FFEF", X"FE19", X"FFA4", X"04AF", X"095B", X"0B16", X"0926", X"0AB3", X"048C", X"0400", X"FE40", X"0142", X"FFCF", X"FFF9", X"FED0", X"FAE8", X"F672", X"F948", X"F8D0", X"FA3F", X"FC63", X"FD1D", X"FD1C", X"FD2C", X"FC62", X"FEC6", X"FF52", X"FF4B", X"00E8", X"FF76", X"048D", X"07A4", X"0C30", X"0890", X"05D6", X"09E9", X"04A9", X"034A", X"FE17", X"0067", X"FF00", X"0015", X"0181", X"FFC4", X"FBCA", X"F95A", X"F954", X"F71D", X"F680", X"F7B7", X"FBF1", X"F9F1", X"FBFE", X"FF3F", X"FFB4", X"0273", X"0090", X"00B1", X"0196", X"0044", X"05E7", X"0287", X"FEAF", X"0557", X"FFBC", X"FF9F", X"00E8", X"FFFC", X"00EB", X"00D5", X"FF43", X"017B", X"01C4", X"FF7F", X"FDE1", X"FC76", X"FCAB", X"FC92", X"FF51", X"01C7", X"04A4", X"002C", X"FFCA", X"FC6E", X"FD09", X"FC8A", X"F9F1", X"F958", X"FD6E", X"FC00", X"FC1E", X"FDB8", X"FE9D", X"0035", X"FE8D", X"00B6", X"0080", X"FE9C", X"0059", X"FEC6", X"FF70", X"FFBC", X"FCE1", X"FC5F", X"FC11", X"FDD7", X"FCD6", X"004F", X"000C", X"FCAD", X"FD2E", X"FF91", X"FDF3", X"FC62", X"FDAB", X"FAD2", X"FDA5", X"FD5F", X"FE2B", X"FE30", X"004D", X"0134", X"00B8", X"FF66"),
        (X"FFC3", X"FFB3", X"FEE8", X"FFE6", X"FF57", X"FFEA", X"0065", X"FF3F", X"00B7", X"00EC", X"FF50", X"0010", X"008B", X"FEA0", X"FFE6", X"004F", X"00DC", X"FF79", X"002F", X"01AA", X"FF99", X"0008", X"FFD1", X"FE3E", X"000B", X"0057", X"00A3", X"FF23", X"FF51", X"00F5", X"FF1C", X"FF6F", X"FF71", X"008B", X"FFEA", X"FEDF", X"FE4C", X"00C3", X"00A3", X"FEE2", X"FCEE", X"FDCF", X"0163", X"0233", X"FC78", X"FCE1", X"01F2", X"0016", X"005C", X"FE34", X"FDC5", X"FE2B", X"0039", X"FF6F", X"FEDC", X"FFED", X"0003", X"FE70", X"00CF", X"FE81", X"FF07", X"0000", X"FF4B", X"FD1E", X"FE2B", X"FB85", X"FBF6", X"F9F4", X"FBB7", X"FFC5", X"00E4", X"FF9E", X"0006", X"FED9", X"01A1", X"02A4", X"0268", X"0053", X"FF95", X"FD5B", X"FC91", X"FD62", X"FFC2", X"FEA5", X"003E", X"FE38", X"FEEB", X"FE0E", X"01F6", X"03B9", X"01EB", X"003D", X"0032", X"00A0", X"004B", X"FF9B", X"FE23", X"FF56", X"FE81", X"0104", X"FED2", X"004C", X"021F", X"FF91", X"01AB", X"0147", X"017A", X"004E", X"FDE2", X"FF08", X"FFB2", X"FF72", X"FF92", X"FF13", X"00F9", X"0263", X"019B", X"0159", X"0160", X"02B3", X"FF3D", X"FF83", X"FF2A", X"FE02", X"FE02", X"FE4F", X"FF63", X"0074", X"FE93", X"FEBC", X"FFF5", X"FF99", X"FFB1", X"0198", X"000F", X"006F", X"03CB", X"02A0", X"FFC0", X"FDC6", X"FEF1", X"00CA", X"0094", X"0362", X"03AB", X"01D5", X"009E", X"0053", X"FDB0", X"FF60", X"FB08", X"FD0C", X"FDB4", X"FE5D", X"FE91", X"FE95", X"FDAC", X"FCCB", X"FE0A", X"FE5F", X"FFEC", X"FE77", X"FF24", X"FFD9", X"02C8", X"038E", X"FFCB", X"FD57", X"01B2", X"0082", X"00FE", X"022B", X"0131", X"0229", X"FEE7", X"FD9C", X"FDEA", X"FE19", X"FE02", X"FD83", X"FC9A", X"FE22", X"FCF1", X"FE5F", X"FE8A", X"FCC1", X"FDC5", X"FDF9", X"FF39", X"FC3E", X"FE17", X"0154", X"050F", X"041F", X"01F7", X"0111", X"FF90", X"01DD", X"FF4C", X"02CF", X"0224", X"013F", X"FE7B", X"FE09", X"FE25", X"FFC3", X"FD42", X"FB6C", X"FC98", X"FA29", X"FA5A", X"FBF1", X"FDBB", X"FD6A", X"FD25", X"FB7F", X"FE22", X"FDB7", X"FD86", X"FFAA", X"00F4", X"0406", X"0252", X"0208", X"FDCB", X"FB42", X"0100", X"02C0", X"012F", X"007B", X"0234", X"018B", X"0081", X"FE84", X"FC39", X"FC03", X"FC6E", X"FE1A", X"FA21", X"FA58", X"FB7C", X"FAD5", X"FF4C", X"FC2D", X"FEDF", X"FEEF", X"FF92", X"FBB8", X"02AA", X"0307", X"02C8", X"029F", X"0011", X"FDDB", X"0097", X"037B", X"00D9", X"FD60", X"024A", X"0251", X"00DC", X"FE05", X"FED8", X"FC92", X"FE64", X"FF50", X"FF0D", X"FF5B", X"FCFB", X"FCFF", X"FD12", X"FDEB", X"00FD", X"01C1", X"0207", X"000C", X"02C3", X"0348", X"03D9", X"FF8C", X"FFC2", X"FEA3", X"FE27", X"03DB", X"0325", X"FE6C", X"0162", X"01F5", X"02CF", X"FF17", X"FEDA", X"FF7C", X"014D", X"056F", X"086B", X"0477", X"0178", X"FF2C", X"0047", X"00A7", X"01DC", X"0202", X"02C8", X"0095", X"0401", X"0582", X"0274", X"FF4B", X"0024", X"FCA2", X"0084", X"058C", X"033D", X"02CC", X"02A0", X"03B2", X"0337", X"0136", X"045E", X"04F9", X"0784", X"0C76", X"0CBB", X"09A9", X"051F", X"04EF", X"03F6", X"0152", X"01D2", X"FF97", X"01A7", X"01F5", X"0344", X"04EA", X"047A", X"0022", X"FFDD", X"FDC6", X"FE76", X"04FF", X"01E8", X"0389", X"051F", X"06C8", X"03B2", X"05AA", X"0627", X"0817", X"0AD5", X"0B55", X"0BC5", X"0A51", X"0883", X"06C0", X"0615", X"037B", X"035A", X"028D", X"0362", X"00C4", X"01FE", X"037C", X"01E4", X"FEDE", X"0144", X"FF9F", X"FE08", X"04BD", X"055F", X"043E", X"07D1", X"0725", X"038C", X"03FF", X"0415", X"0787", X"0790", X"074E", X"0773", X"08A3", X"0694", X"08FC", X"084B", X"05D2", X"04BF", X"0368", X"0211", X"0124", X"0044", X"0016", X"FD8D", X"FE9D", X"FDE5", X"0210", X"00EE", X"06E2", X"067F", X"04AA", X"06A8", X"0265", X"01D9", X"0128", X"0310", X"0493", X"0636", X"02FA", X"03BB", X"04CC", X"072F", X"0710", X"085E", X"089E", X"051C", X"03A8", X"027D", X"024E", X"026B", X"0065", X"F99E", X"FDCC", X"FEFB", X"02BA", X"0411", X"0562", X"04BC", X"003C", X"0180", X"0016", X"FD80", X"FF78", X"0157", X"042A", X"03B2", X"0329", X"02B2", X"0359", X"03AA", X"055C", X"0739", X"0828", X"024F", X"0010", X"028D", X"0234", X"FF89", X"FCDA", X"F938", X"FD2E", X"0141", X"0286", X"02D8", X"061C", X"001F", X"FB87", X"FD9A", X"FFA3", X"FF81", X"00A0", X"004C", X"0226", X"036D", X"0153", X"048D", X"030E", X"02DC", X"05BD", X"034A", X"0327", X"FDE0", X"FEA2", X"00DD", X"011D", X"000D", X"F96E", X"FA47", X"FD40", X"000A", X"01E7", X"04BE", X"039B", X"FDC5", X"FCA3", X"FF69", X"FFB1", X"00D3", X"FF2D", X"FF01", X"FFBC", X"02CC", X"02DF", X"02D3", X"0428", X"0532", X"02C4", X"0068", X"028E", X"FF32", X"FE21", X"011B", X"024D", X"FECE", X"F91B", X"F9EC", X"FDB1", X"FF3F", X"0084", X"03D3", X"045F", X"FC92", X"FE76", X"FF13", X"FEFF", X"FFAF", X"FEB9", X"FF12", X"FEF8", X"FF33", X"00DB", X"028C", X"0391", X"023F", X"FEE1", X"FDD5", X"FF2C", X"FF0B", X"FE35", X"FFE0", X"FF6D", X"FB82", X"F9D4", X"FAF9", X"FEAA", X"FFF6", X"0022", X"00FF", X"0269", X"FD90", X"0185", X"FD01", X"FD01", X"FEB4", X"FE8E", X"FE4F", X"FC60", X"FB7A", X"FD88", X"FFFF", X"019A", X"0116", X"FE4D", X"FF41", X"0065", X"FD38", X"FF53", X"FF27", X"0175", X"FE13", X"F95C", X"FC46", X"FF61", X"FEDE", X"0108", X"FF1D", X"0047", X"FAB0", X"FC57", X"FCCB", X"FDC2", X"FDB1", X"FBE8", X"FC88", X"FAF4", X"FA1D", X"FBB4", X"0038", X"0139", X"FD1A", X"FDC3", X"FEB9", X"FDC7", X"FC60", X"FE28", X"FE25", X"FC88", X"FBD3", X"FAF7", X"FD27", X"012D", X"0052", X"FF55", X"FFF3", X"FF9C", X"FC7B", X"FC7B", X"FED8", X"FEA7", X"FD17", X"FC55", X"FC71", X"F8E6", X"F96C", X"FCE9", X"FF8F", X"FEC7", X"FE0D", X"FC17", X"FE0C", X"FADA", X"FC4F", X"FCDF", X"FCED", X"FA40", X"FA87", X"FBE7", X"FCC3", X"0121", X"018C", X"FF0C", X"FE48", X"004D", X"FF0B", X"FC4C", X"FDD5", X"FDF5", X"FD56", X"FC2F", X"FD39", X"FBD3", X"FC29", X"FD1E", X"FEEA", X"0057", X"FE4C", X"FF1A", X"FE81", X"FC2C", X"FAD5", X"FA98", X"FB85", X"FCE7", X"FB0C", X"FCEA", X"01C6", X"FECF", X"FEC9", X"FF93", X"02B3", X"04AB", X"0227", X"010D", X"FF5D", X"FFA4", X"0235", X"FF2E", X"FF73", X"FC28", X"FC0E", X"FE88", X"FE74", X"00C2", X"024B", X"011B", X"FE54", X"FE01", X"FC73", X"FA50", X"FBF5", X"FE4B", X"FE04", X"FD2B", X"018A", X"FF61", X"FE67", X"FE36", X"FFCA", X"06DD", X"0391", X"0039", X"037F", X"02E1", X"0242", X"01D6", X"0161", X"01B0", X"FE8A", X"FFA8", X"0150", X"FEF3", X"012E", X"FE52", X"FE68", X"0064", X"004A", X"FF1E", X"FEA4", X"0088", X"FA2E", X"FB4E", X"FE94", X"FFCC", X"0114", X"000F", X"0129", X"FE0A", X"FE46", X"0010", X"01F4", X"FD4D", X"FEEF", X"00A4", X"028E", X"00DE", X"0059", X"0275", X"0368", X"030D", X"0344", X"0398", X"0644", X"0791", X"04A7", X"001D", X"0119", X"03E5", X"FE4E", X"FE2C", X"FF4E", X"FF4A", X"00D3", X"FFC8", X"0121", X"FF77", X"0095", X"010D", X"FF0F", X"FCDE", X"F844", X"F7AA", X"F762", X"FA91", X"FC82", X"FCEC", X"FBE5", X"FAC5", X"FCD3", X"FF7F", X"0004", X"01C9", X"0313", X"047A", X"0202", X"0126", X"FF50", X"007D", X"FFF8", X"002E", X"0051", X"FF94", X"019E", X"FF99", X"FF31", X"0033", X"FEA1", X"FD07", X"FCC6", X"FBCF", X"FE2E", X"FDE1", X"FC02", X"F9AB", X"F8AC", X"F9CA", X"F98C", X"F9D5", X"FDBE", X"FE36", X"FF6F", X"00C3", X"01EE", X"FDC4", X"FFDE", X"FF70", X"FFF0", X"0035"),
        (X"FF31", X"01CD", X"FFCA", X"FF80", X"0037", X"0021", X"0045", X"00E3", X"0094", X"0034", X"002A", X"FF5B", X"FF90", X"FF4E", X"FE48", X"FE65", X"0154", X"0036", X"FF7D", X"FFC8", X"00DC", X"0026", X"00A7", X"0124", X"00EA", X"000F", X"017F", X"FF17", X"FE47", X"006B", X"0005", X"FF31", X"FF4F", X"FFD1", X"00DA", X"FFEB", X"029E", X"024B", X"0377", X"0268", X"0361", X"01F6", X"FEFE", X"FDC3", X"FC75", X"011C", X"0179", X"039C", X"04DA", X"0139", X"0372", X"008D", X"FF82", X"0078", X"FE11", X"FFF9", X"00B0", X"00FE", X"00B1", X"FFD7", X"FFBA", X"018D", X"FF59", X"0080", X"00D0", X"008E", X"00DE", X"0460", X"0098", X"0123", X"0117", X"FE41", X"FDE8", X"0273", X"041E", X"03DA", X"05B9", X"06CB", X"070B", X"0226", X"0231", X"FFAB", X"FE12", X"0042", X"FF74", X"001D", X"FF3A", X"FEDA", X"00F6", X"04E1", X"033E", X"061E", X"03B0", X"01FF", X"039A", X"033F", X"017A", X"FE8B", X"0177", X"01E0", X"0531", X"0443", X"0694", X"07DE", X"08B4", X"07C8", X"079C", X"083A", X"05FA", X"FCC3", X"FE32", X"FFC7", X"009D", X"0071", X"FD69", X"00D2", X"0419", X"05E9", X"04EB", X"06EE", X"03DB", X"01D1", X"FFD3", X"0086", X"FD2E", X"FD77", X"FD3A", X"006B", X"050F", X"05DA", X"06DD", X"0776", X"067E", X"07CA", X"07B9", X"0541", X"027F", X"FFFB", X"0255", X"0274", X"00EC", X"0111", X"FDB6", X"FF27", X"0460", X"07CE", X"0792", X"051C", X"06C7", X"0451", X"018B", X"00EB", X"01E7", X"01E5", X"FFDD", X"0141", X"04B1", X"07CD", X"0769", X"073C", X"05B3", X"0356", X"0162", X"0019", X"004E", X"02DC", X"FF44", X"FFFE", X"FFEC", X"0075", X"02B5", X"FFDB", X"03AB", X"0A7E", X"0900", X"094B", X"0987", X"07BA", X"038A", X"0291", X"02E5", X"04FD", X"037F", X"0535", X"071F", X"0819", X"04B3", X"05C9", X"02F7", X"030B", X"0107", X"FD0A", X"0063", X"00AD", X"FD07", X"FF6F", X"00CD", X"01CB", X"FFEE", X"0343", X"0698", X"09CD", X"0B63", X"0C9B", X"0D83", X"0B00", X"05C0", X"02FE", X"016B", X"043D", X"01DB", X"0435", X"054E", X"04D7", X"02FE", X"023C", X"01E6", X"0115", X"FEB0", X"FCCA", X"FE43", X"FE51", X"FDF8", X"FE9B", X"FF6F", X"FF2B", X"005E", X"0422", X"07E5", X"0611", X"064D", X"08E6", X"0885", X"091A", X"0406", X"0035", X"01BE", X"FEEB", X"FF00", X"FF03", X"0067", X"FE20", X"FFDB", X"FFEC", X"00EC", X"FF29", X"FD71", X"FCAA", X"FC03", X"FCF0", X"FF0E", X"FDEB", X"00B7", X"0117", X"FDC8", X"0488", X"06E6", X"0787", X"038B", X"047F", X"052D", X"0515", X"FF6C", X"FF04", X"FE6C", X"FC96", X"F7FC", X"F54C", X"F996", X"FB06", X"FE4F", X"00AA", X"0253", X"FFF1", X"0032", X"001B", X"FCA2", X"FAB1", X"FB94", X"FBEB", X"FF82", X"FE6D", X"FE86", X"055A", X"06D7", X"04B5", X"041F", X"007E", X"02D8", X"01A6", X"FF4A", X"FC84", X"FC7C", X"FA79", X"F73E", X"F5E9", X"F6EF", X"FC39", X"025C", X"0326", X"02E3", X"027D", X"00C8", X"FFA3", X"F8A6", X"F473", X"F72A", X"FF6A", X"0066", X"0008", X"01D6", X"0525", X"03AC", X"01F8", X"0395", X"0224", X"034C", X"0472", X"03B9", X"FDAE", X"FD45", X"FCA6", X"F9AD", X"F99B", X"FA55", X"006A", X"0449", X"03F6", X"0359", X"012E", X"FFF5", X"FE26", X"FCE9", X"F5B4", X"FA28", X"FFFC", X"FF4F", X"FFE9", X"0330", X"0461", X"01CF", X"0537", X"04B4", X"05E7", X"0420", X"0395", X"033A", X"0247", X"0057", X"FF54", X"FCCE", X"F927", X"FFA6", X"02A4", X"048C", X"04BF", X"05A9", X"0589", X"0618", X"0678", X"0419", X"FDBB", X"F9AF", X"FC88", X"0106", X"00C9", X"0223", X"017A", X"025B", X"0532", X"057D", X"03E5", X"FF4F", X"FF86", X"009D", X"FFC5", X"01AE", X"FF83", X"FC47", X"FDA0", X"FF99", X"026F", X"068B", X"0AB1", X"0A63", X"087A", X"0583", X"051F", X"00EF", X"FCEF", X"F67D", X"FDDF", X"FFF5", X"00B9", X"FF3A", X"FEE1", X"0222", X"021E", X"03BC", X"01C5", X"FC9C", X"FCCF", X"FF0A", X"026F", X"02BE", X"0098", X"FDC6", X"FE9A", X"FE63", X"030D", X"0823", X"0A67", X"082F", X"067D", X"0070", X"FEDB", X"FBD7", X"FD23", X"F782", X"FC84", X"0021", X"FEE6", X"FFBC", X"FFA0", X"0247", X"001D", X"00EC", X"FF33", X"FCDF", X"FD4D", X"FE4A", X"004E", X"006F", X"FEC6", X"FDFF", X"FD22", X"FD25", X"04EE", X"07D1", X"0906", X"085E", X"02A6", X"FF09", X"FE09", X"FA83", X"F9A3", X"F7AD", X"FE4A", X"0017", X"0163", X"00E0", X"0001", X"011F", X"FEB7", X"FFD5", X"FFCC", X"FD9A", X"FE57", X"FF0A", X"FFE3", X"0038", X"FD2D", X"FBE6", X"FD4D", X"024E", X"0589", X"06A1", X"0784", X"033F", X"FEFC", X"FB32", X"FA24", X"FA72", X"F966", X"F5D9", X"FC05", X"0124", X"FF3B", X"02D7", X"FEDA", X"FFEC", X"FCC3", X"FB66", X"FD36", X"FD98", X"FDB3", X"FD64", X"FF84", X"FCFC", X"FCCD", X"FC33", X"FED7", X"022B", X"06D6", X"03A3", X"0328", X"0062", X"FF14", X"FC20", X"FB68", X"F993", X"FB54", X"F98E", X"FA91", X"00B2", X"014D", X"026C", X"FF32", X"FE61", X"FCE0", X"FDF5", X"FCE6", X"FE5D", X"FD72", X"FDE3", X"0033", X"FB3A", X"F9A5", X"FC01", X"0033", X"0428", X"027F", X"0158", X"0240", X"FEEB", X"FD7F", X"FB1F", X"FA55", X"F843", X"FAB9", X"FE01", X"FD2A", X"FF71", X"FF87", X"01B3", X"FEAB", X"0072", X"0003", X"FF35", X"FF6E", X"FD7E", X"FD8B", X"FE40", X"FC99", X"FD38", X"FB0D", X"FC8D", X"011B", X"0192", X"0011", X"0293", X"FFDC", X"FE82", X"FD79", X"FD9F", X"F9A2", X"FA19", X"F8CA", X"FC72", X"FC36", X"0052", X"0106", X"03F5", X"02C9", X"FFC3", X"049B", X"FFBB", X"FE8A", X"FC06", X"FD6E", X"FFF2", X"FBA5", X"0031", X"00B6", X"0245", X"016B", X"0002", X"0116", X"FF6C", X"FDF7", X"FF19", X"FD04", X"FC67", X"FE55", X"FB13", X"FC14", X"FE07", X"FF73", X"FF25", X"FED0", X"0312", X"01EF", X"FD71", X"FF9F", X"FF45", X"FF56", X"0088", X"FEF5", X"FF27", X"041A", X"042B", X"05DE", X"0558", X"0229", X"03B3", X"FEF8", X"FD17", X"FE95", X"FCE8", X"FCBF", X"FFCC", X"FF1D", X"FBD8", X"FB06", X"FE9E", X"00BA", X"FFF6", X"FFBB", X"02F6", X"025F", X"FCFC", X"FD6F", X"FFEC", X"01E3", X"01C0", X"0050", X"028C", X"0516", X"06D2", X"06DE", X"0541", X"038C", X"021C", X"FD9F", X"FAF3", X"FC0F", X"FBE5", X"FC68", X"0028", X"FC98", X"FC5F", X"FA27", X"FD53", X"FFE1", X"0014", X"0056", X"FFF9", X"03C3", X"FFE2", X"FD40", X"FFB4", X"006D", X"0264", X"033B", X"0380", X"0398", X"0410", X"0687", X"0692", X"028F", X"FFD5", X"FD75", X"FDA9", X"FEEE", X"FE80", X"0017", X"FE61", X"FE3F", X"FB2E", X"FB41", X"FDC3", X"FF73", X"010B", X"FF8D", X"00EF", X"047D", X"0375", X"017D", X"0488", X"06F4", X"0611", X"0674", X"0580", X"072D", X"06AC", X"07F6", X"063F", X"0622", X"07DB", X"0110", X"017D", X"028F", X"04F6", X"FEF0", X"FDDA", X"FF8D", X"FD20", X"FDB2", X"FDE0", X"FEB1", X"FEAB", X"FFD1", X"0037", X"022F", X"067E", X"0760", X"0900", X"0957", X"087F", X"06E8", X"0790", X"0731", X"0750", X"05F5", X"056F", X"0748", X"0A19", X"0622", X"04CD", X"076A", X"03E8", X"02CC", X"0320", X"FECE", X"FD98", X"FD64", X"FD18", X"0119", X"014C", X"FE58", X"FF83", X"00E0", X"02D2", X"04C2", X"0894", X"0756", X"083F", X"08AE", X"07EA", X"0493", X"02B0", X"03B8", X"03C4", X"05B0", X"034C", X"03AE", X"0536", X"0629", X"04A9", X"0351", X"021B", X"0176", X"008F", X"0008", X"FFAF", X"FF54", X"015A", X"FFE0", X"005D", X"FFCC", X"FFD9", X"015A", X"0262", X"01B3", X"046D", X"00BD", X"FF93", X"FE66", X"000F", X"019C", X"0531", X"01FD", X"01B5", X"03A9", X"0259", X"0197", X"008E", X"01A8", X"022D", X"FFDC", X"FEFE", X"FFC5", X"FF1D", X"FF9C"),
        (X"0147", X"FFF3", X"FF49", X"00B2", X"FFE6", X"FF81", X"FFB8", X"FFA2", X"FED3", X"007A", X"0116", X"FFC9", X"FE90", X"00D5", X"0094", X"FF39", X"0011", X"00B4", X"FEF7", X"FFA7", X"FFBB", X"FE9E", X"01A2", X"0076", X"0137", X"FFD9", X"01DC", X"00C9", X"FEF6", X"003F", X"0042", X"FF98", X"FFED", X"0120", X"FE36", X"FDB5", X"FB83", X"FACE", X"FC34", X"F9D2", X"F8F0", X"FCF8", X"0030", X"012B", X"FD70", X"FB82", X"FB2C", X"FA96", X"FB42", X"FE4E", X"FC65", X"FD20", X"0050", X"0001", X"FFFB", X"FFB9", X"FF0E", X"FFEF", X"FFA9", X"FE34", X"FE2F", X"FF9A", X"FFCF", X"FE4B", X"FC11", X"FB06", X"FA04", X"F885", X"F906", X"FA7F", X"FB95", X"FF88", X"FE89", X"FBFD", X"FAB8", X"F629", X"F56C", X"F767", X"F65F", X"FBC0", X"FE79", X"007E", X"FEF7", X"0084", X"FFDA", X"FFF4", X"0200", X"FE94", X"FEEA", X"FF1C", X"FDA6", X"FCA9", X"FD79", X"FDC6", X"FBAB", X"FA12", X"FC89", X"FA84", X"F82B", X"FBB8", X"FB66", X"FB13", X"FB60", X"F8EE", X"F6D5", X"FA81", X"FD22", X"FF62", X"FC16", X"FD5D", X"00CC", X"FECC", X"FE74", X"0070", X"0053", X"FE33", X"FCBF", X"FEA6", X"FEC5", X"FF56", X"006D", X"FF7F", X"FEF8", X"FE3D", X"FFEE", X"FFA8", X"FFB6", X"001F", X"0062", X"0191", X"FF85", X"00C6", X"0243", X"00A1", X"FD2B", X"FE92", X"FF32", X"FF87", X"03BF", X"017A", X"FDB0", X"FFB1", X"FED6", X"FEC6", X"FF19", X"FFFC", X"FF91", X"FEBE", X"FEFF", X"FF71", X"FF40", X"FF2A", X"0094", X"008B", X"020F", X"FF32", X"FF18", X"FF54", X"00B8", X"0107", X"027B", X"02EE", X"00AC", X"0158", X"00CE", X"0196", X"006F", X"02A4", X"FE69", X"005B", X"0296", X"00FB", X"FF92", X"0120", X"FFE8", X"0051", X"012B", X"0230", X"FF75", X"FF27", X"002C", X"FD61", X"FBF9", X"FD30", X"FBB3", X"FC9C", X"FDCF", X"FF1E", X"FF8E", X"0348", X"0319", X"037D", X"0161", X"003B", X"FEFF", X"01AB", X"FFC4", X"005B", X"0514", X"0449", X"042E", X"001B", X"0468", X"0319", X"02CB", X"00F0", X"02D2", X"00B5", X"FF78", X"FE47", X"FBCE", X"FB72", X"FB74", X"FDEC", X"FF1A", X"FF59", X"0158", X"02D8", X"04AB", X"033B", X"03D3", X"FFBA", X"FDB7", X"013E", X"FE4E", X"0248", X"0796", X"0430", X"052D", X"04BB", X"04BE", X"06EE", X"04E2", X"02EB", X"0334", X"0348", X"0320", X"019C", X"FE92", X"FEEC", X"FE02", X"0014", X"FF47", X"0216", X"0102", X"0217", X"0328", X"05DE", X"050B", X"FFCA", X"01DF", X"0230", X"01B1", X"02A9", X"032E", X"024E", X"07B7", X"08F5", X"0704", X"049B", X"0477", X"03F8", X"0482", X"057F", X"0268", X"000E", X"0067", X"000D", X"02D4", X"00D2", X"00FD", X"02AE", X"01F6", X"0314", X"050B", X"04E1", X"0310", X"0140", X"0263", X"FDD5", X"005C", X"055A", X"059B", X"04A7", X"062D", X"0608", X"0704", X"0540", X"02A8", X"0331", X"02EC", X"01BF", X"0084", X"00A6", X"0224", X"02AF", X"01C7", X"0132", X"00B5", X"006B", X"0065", X"00B4", X"01F0", X"03CD", X"0026", X"FE1D", X"0058", X"0215", X"022E", X"0469", X"06A3", X"0320", X"036D", X"0317", X"0183", X"048E", X"03B3", X"01AB", X"FD96", X"FB69", X"F983", X"FD37", X"014A", X"FF79", X"FD67", X"FAAD", X"FBEB", X"FEA8", X"FDAA", X"FDF8", X"0099", X"FECD", X"00C4", X"0244", X"04FF", X"00D4", X"011C", X"032A", X"04B5", X"0045", X"FF14", X"FDE3", X"FD9E", X"FEAF", X"FDFA", X"FC1C", X"F6B1", X"F6E0", X"F8A9", X"FD11", X"FE16", X"FDE0", X"FB25", X"F949", X"FBC0", X"FCE2", X"FF4B", X"01A9", X"FF84", X"FF50", X"0421", X"0820", X"08C1", X"0438", X"012D", X"03D1", X"04F1", X"FB44", X"F882", X"F78E", X"F790", X"F7C4", X"F896", X"F857", X"F623", X"F859", X"FB95", X"FF83", X"FF5B", X"0061", X"FAB8", X"FBF9", X"FDB2", X"FE45", X"FE44", X"FE76", X"FE3F", X"FEDA", X"FF10", X"074A", X"08A9", X"04FC", X"017B", X"FDAC", X"0004", X"F9D4", X"F3D1", X"F1D0", X"F337", X"F363", X"F2C6", X"F64F", X"F8C7", X"FC36", X"FFD4", X"04F2", X"01E4", X"0044", X"FE9C", X"FE9A", X"FEA5", X"FE04", X"FCA9", X"FC1E", X"FD19", X"FA25", X"FBB7", X"04D0", X"09F4", X"0561", X"FFB0", X"FCBB", X"FDA8", X"FA9E", X"F6B1", X"F1E5", X"F2B1", X"F294", X"F537", X"FA10", X"FD25", X"00F0", X"049F", X"0656", X"059E", X"007F", X"01AD", X"FFF6", X"FF7F", X"FE3A", X"F813", X"F9D2", X"FA30", X"FBB6", X"FD6F", X"060C", X"09EF", X"03CC", X"0081", X"FCF0", X"FA9D", X"FCD2", X"F6D2", X"F568", X"F841", X"F8CE", X"FC49", X"FF1E", X"0184", X"02C6", X"04C6", X"06EA", X"04F9", X"04FA", X"04BC", X"0086", X"FE8F", X"FC40", X"FAC0", X"FB4B", X"FAA6", X"FD4E", X"FDAA", X"0651", X"0A00", X"0574", X"FFA3", X"FD9E", X"FC29", X"FD01", X"FAD8", X"FB19", X"FBB9", X"0001", X"FFD6", X"01AB", X"01F2", X"0222", X"0446", X"05C5", X"0511", X"03C2", X"01AE", X"FEC9", X"FE2C", X"FDC1", X"FDB8", X"FD3D", X"FC44", X"FD62", X"0113", X"0778", X"0743", X"039D", X"000A", X"FF84", X"FCF2", X"FF18", X"FC35", X"FDFE", X"0080", X"01AF", X"0236", X"0337", X"02EF", X"0299", X"0566", X"0687", X"045A", X"0223", X"FE5B", X"FE5C", X"FE4E", X"FD9D", X"FF59", X"FB80", X"FC67", X"FD50", X"0363", X"054A", X"0527", X"01B2", X"FFC2", X"FE5E", X"FB00", X"FE76", X"FEA6", X"FF38", X"0223", X"038A", X"0362", X"064F", X"04CC", X"04F8", X"043B", X"0501", X"0187", X"006B", X"FE27", X"FED4", X"FF11", X"FE46", X"FE30", X"FE93", X"FD61", X"01AF", X"0300", X"06BE", X"077A", X"02E9", X"0062", X"FCE0", X"FCCF", X"FD00", X"FBAC", X"FDB2", X"01FD", X"0415", X"03A9", X"047E", X"04E0", X"043D", X"0307", X"023B", X"0047", X"FF1B", X"FE2E", X"FEF6", X"FECD", X"00A2", X"FE96", X"FF66", X"FFA0", X"024E", X"02B1", X"008C", X"052D", X"004B", X"0087", X"0004", X"FE63", X"FEF9", X"FC82", X"FE54", X"028E", X"022E", X"0219", X"02F6", X"00DA", X"0175", X"FF53", X"FF69", X"FEFA", X"FE37", X"FEF6", X"0194", X"0057", X"0210", X"01BF", X"00AC", X"0209", X"0353", X"022A", X"0233", X"01F5", X"FFF1", X"0015", X"FF07", X"FE03", X"FBA8", X"005A", X"013B", X"02FE", X"01E0", X"0087", X"0138", X"FF9E", X"00B8", X"FFE1", X"FFCB", X"01B8", X"009D", X"003B", X"0050", X"01AD", X"014C", X"00EF", X"0288", X"0285", X"010B", X"0066", X"01A5", X"FCCD", X"FEA3", X"FF75", X"FF2D", X"FCA6", X"F7D4", X"FAE6", X"FC41", X"FCD6", X"FDC5", X"FDB1", X"0013", X"FE09", X"0074", X"0280", X"0271", X"0314", X"0309", X"02A2", X"012F", X"01EA", X"0231", X"023C", X"029E", X"00FA", X"FD9D", X"FDB5", X"0051", X"FDC8", X"0020", X"FFA8", X"010D", X"FDAD", X"F849", X"F4E9", X"F6BE", X"FA16", X"F825", X"FA13", X"FC15", X"FC73", X"0015", X"0174", X"00A6", X"0315", X"01C9", X"00C0", X"FECB", X"004A", X"01B5", X"0081", X"FE3D", X"F9E3", X"F95D", X"01E7", X"036A", X"0182", X"FFBC", X"FFCF", X"00C9", X"FD33", X"018B", X"FA30", X"F7C7", X"F983", X"F8FC", X"F893", X"FA1C", X"FB96", X"FD31", X"FBBC", X"FC92", X"FEEE", X"FFC7", X"FE87", X"FE3D", X"FBC2", X"FA65", X"F9D1", X"FB5D", X"F827", X"F979", X"FB6C", X"FE4D", X"0294", X"FF45", X"00D1", X"FFD0", X"0039", X"FDD6", X"FCA3", X"F9EA", X"FAE7", X"FBAE", X"0040", X"FDF6", X"FC42", X"FE7E", X"FC02", X"FA20", X"F901", X"FB26", X"F9B7", X"F981", X"F9C3", X"F8EF", X"F8BD", X"FC75", X"FFE0", X"FFE0", X"FF42", X"012E", X"01D2", X"01C6", X"0070", X"0019", X"00C5", X"FFB4", X"014D", X"026C", X"00F5", X"010B", X"01BC", X"02F6", X"01FF", X"01F4", X"009F", X"099A", X"039A", X"0618", X"08B8", X"0755", X"02B7", X"026C", X"FEB1", X"FEE7", X"FFA8", X"0150", X"FEFF", X"01B1", X"FFFF", X"004C"),
        (X"0045", X"FF8F", X"FFCF", X"FF54", X"0071", X"00DD", X"FED3", X"FF9B", X"014D", X"FF6D", X"FF58", X"0032", X"000B", X"00EA", X"0225", X"00C6", X"005D", X"FF34", X"012D", X"0123", X"FF2C", X"006E", X"FFB5", X"FF7F", X"FFAA", X"FE99", X"0074", X"FF54", X"007B", X"FF0A", X"0170", X"00C3", X"0078", X"00DF", X"FF47", X"FEA6", X"FDEE", X"FC92", X"FCF8", X"0096", X"FE5E", X"00A5", X"00ED", X"0309", X"034C", X"FFF6", X"008A", X"FD31", X"FD9F", X"0084", X"FEBD", X"FFBB", X"FFD0", X"00C9", X"000E", X"FE39", X"FFE3", X"FF67", X"FF28", X"0054", X"FFC5", X"0023", X"FEBA", X"FECB", X"FF31", X"00F8", X"0288", X"011F", X"010A", X"022A", X"00D0", X"016F", X"0328", X"FED4", X"FB4F", X"FAA8", X"FB01", X"FC28", X"FC26", X"FF58", X"032F", X"028B", X"FFA9", X"FE53", X"FF52", X"FF77", X"03EE", X"006A", X"FE6C", X"00DE", X"FF3D", X"0103", X"0258", X"01F1", X"0219", X"0383", X"041A", X"0412", X"02DD", X"FED4", X"FEBA", X"FC2B", X"F8B9", X"F640", X"F763", X"F9AE", X"F743", X"FCB8", X"FF48", X"010E", X"FF84", X"FF8F", X"004C", X"FF1F", X"02FC", X"000F", X"FFD0", X"0079", X"02DD", X"034E", X"0508", X"067A", X"06F3", X"0514", X"032A", X"01AD", X"02A6", X"012B", X"FCF2", X"FAAE", X"FC55", X"F768", X"F8C3", X"F7B3", X"F7EF", X"F900", X"F978", X"FDAF", X"FEC2", X"FDC6", X"012F", X"FF96", X"0293", X"00AB", X"01D7", X"FF9B", X"FEB5", X"FDAD", X"0045", X"01C4", X"03B6", X"05EF", X"0396", X"0408", X"0151", X"0172", X"FEAE", X"FFF0", X"FFA5", X"004E", X"00E4", X"FE6B", X"FCAD", X"F98D", X"FB28", X"FDF9", X"FD65", X"FCE0", X"FFA3", X"0050", X"FDFC", X"FE70", X"FE22", X"F9BC", X"FD57", X"FB4B", X"FE16", X"00BB", X"06A5", X"08C8", X"0815", X"0803", X"061B", X"06DB", X"06F0", X"0795", X"0993", X"063D", X"0802", X"04CA", X"FEBB", X"FB12", X"F895", X"FE90", X"FE9E", X"FE42", X"0003", X"FE38", X"FCC9", X"FBA3", X"FCE6", X"F8A5", X"F8AF", X"F8C1", X"FCBD", X"FF78", X"04AC", X"0798", X"0BEE", X"0BC6", X"0BED", X"0AA9", X"0B63", X"0B3D", X"09A9", X"0A70", X"07C8", X"060C", X"FFDD", X"FC46", X"F896", X"FC8C", X"FD71", X"FFCB", X"0006", X"FE66", X"FCFC", X"F965", X"FB73", X"FA1A", X"FA37", X"F9EC", X"FB93", X"FFB8", X"008B", X"035A", X"0522", X"096C", X"0A70", X"0AB3", X"09F3", X"06D7", X"0627", X"0629", X"020A", X"01F2", X"0149", X"FC93", X"FAB2", X"FB3A", X"FFEB", X"016E", X"FE1E", X"FBBD", X"FAFE", X"FB9D", X"FAB7", X"FC04", X"FD1D", X"FD68", X"FCE8", X"FCA2", X"FEAB", X"FCAB", X"FE3A", X"0118", X"0498", X"0439", X"FFCB", X"028C", X"FF61", X"0069", X"FDD7", X"FD16", X"FFAF", X"FD39", X"FB9C", X"FB14", X"FD6E", X"FD91", X"FF7C", X"FC8A", X"F966", X"FCD5", X"FB61", X"FF48", X"00E5", X"FD36", X"FE41", X"FB35", X"FCD9", X"FC07", X"FB09", X"FA88", X"FDB1", X"FB65", X"FA94", X"FE84", X"FFD9", X"FEA4", X"FE80", X"FE04", X"FED6", X"0194", X"FD03", X"FBB6", X"FD71", X"FF67", X"FEE5", X"FBE9", X"F92C", X"FB4E", X"FD33", X"0319", X"012A", X"0054", X"FE6F", X"F9FF", X"FAE9", X"FB28", X"F887", X"FC1E", X"0139", X"FD12", X"FC6D", X"0100", X"009C", X"0017", X"0279", X"01E7", X"024B", X"01DE", X"03B5", X"00B3", X"0272", X"007D", X"FD9C", X"FE02", X"F89E", X"FCDE", X"0019", X"022C", X"FFEF", X"FFF3", X"FEFB", X"FD0D", X"FB65", X"F8D3", X"F736", X"FF93", X"0392", X"FFAC", X"FE74", X"013E", X"02F2", X"029F", X"025F", X"01F6", X"01CD", X"01EE", X"01F3", X"030E", X"020C", X"FF29", X"FF38", X"FEDC", X"FAC9", X"0058", X"02E3", X"0031", X"FDA9", X"FDE2", X"FCBA", X"FDF9", X"FB4C", X"F8F6", X"F909", X"02C0", X"04A5", X"006C", X"FE24", X"FEDC", X"0006", X"0083", X"0086", X"FF02", X"FF11", X"FD14", X"FB09", X"011D", X"0325", X"0147", X"FEBD", X"FEA0", X"FD63", X"FEFC", X"01D6", X"FC7E", X"FD86", X"FF30", X"FE54", X"FD58", X"FC16", X"F9E8", X"FCFB", X"02C4", X"029E", X"0060", X"FD6C", X"FC21", X"FE70", X"FDF2", X"FD53", X"FDDC", X"FC13", X"FBE5", X"F9F8", X"FEAE", X"069A", X"019A", X"FEDE", X"FF50", X"FC10", X"FE20", X"0199", X"0006", X"FC68", X"FDE6", X"FE94", X"FDF6", X"FEAC", X"FBB9", X"FF27", X"013C", X"0127", X"FD56", X"FBDD", X"FC5B", X"FE94", X"FD8B", X"FB94", X"F944", X"F9EB", X"FAB0", X"FE7B", X"FE14", X"0382", X"020F", X"006A", X"FF74", X"015C", X"028D", X"056F", X"0162", X"FF29", X"FE9D", X"FFCC", X"FEFD", X"FF0D", X"FE9D", X"FF55", X"FF79", X"FEEC", X"FCFB", X"FD7D", X"FC2A", X"FBA4", X"FB4C", X"FA19", X"F940", X"FC37", X"FC81", X"FCCD", X"01A6", X"0391", X"03CB", X"FF77", X"004C", X"0155", X"05A3", X"03B7", X"002A", X"FF86", X"FD9E", X"0128", X"FE1B", X"FF44", X"0013", X"00B1", X"001C", X"FC5D", X"FDC1", X"FE29", X"FE51", X"FAA0", X"FD91", X"FD88", X"FBBE", X"00BE", X"FDFE", X"0031", X"0327", X"0540", X"0140", X"0143", X"FF98", X"01DB", X"0514", X"019B", X"0013", X"009A", X"FDDD", X"FE9E", X"FDB3", X"FF5D", X"FEBF", X"FC46", X"FE2B", X"FD91", X"FDE4", X"FFCB", X"FF94", X"007F", X"0247", X"01B7", X"0200", X"03E8", X"0425", X"02B9", X"04DE", X"0446", X"017B", X"FFE1", X"FD77", X"0230", X"0389", X"02C7", X"026F", X"01CF", X"0270", X"008B", X"FF77", X"FD79", X"FAF6", X"FCE9", X"FD7B", X"FDEA", X"FE22", X"FF01", X"FFDB", X"0208", X"02A1", X"02CD", X"039D", X"076B", X"04D2", X"04BE", X"073B", X"0442", X"0057", X"00B1", X"FBA3", X"0268", X"037D", X"058A", X"07F1", X"050C", X"05DD", X"03F1", X"0104", X"FEE4", X"FCEB", X"FD8B", X"FEF0", X"FDC1", X"FE4B", X"FEB3", X"FF44", X"001F", X"02A1", X"0526", X"0658", X"0824", X"0598", X"0704", X"0609", X"03DE", X"00A1", X"0034", X"0137", X"02A6", X"058F", X"0891", X"0814", X"0A0B", X"09E3", X"0274", X"038B", X"0046", X"FE70", X"FBC7", X"FD83", X"FEEF", X"FE5A", X"FFB9", X"FF58", X"0136", X"0373", X"04C6", X"059A", X"0678", X"06F0", X"0609", X"0398", X"FD23", X"FFA7", X"018F", X"0027", X"021E", X"03BF", X"05C0", X"093F", X"0902", X"0839", X"063D", X"04DA", X"0235", X"00BE", X"00F0", X"00C0", X"016B", X"FF3F", X"FE86", X"01B3", X"0328", X"00BB", X"042C", X"0311", X"062E", X"069B", X"04FB", X"0272", X"FCA9", X"0101", X"00DA", X"FFB6", X"01F5", X"0414", X"0322", X"03CD", X"03DF", X"03C8", X"058A", X"0364", X"03B4", X"03A1", X"06D5", X"04BC", X"0298", X"033D", X"03E1", X"0223", X"01E9", X"049A", X"011B", X"01F2", X"0462", X"0417", X"0549", X"0073", X"FE55", X"FFC5", X"0116", X"00B2", X"006A", X"00D6", X"017C", X"FFAD", X"FDE6", X"027D", X"0386", X"0235", X"0328", X"0435", X"04C1", X"05CA", X"0254", X"0365", X"025C", X"0303", X"02A5", X"0138", X"03B6", X"0404", X"036D", X"03AE", X"0298", X"0185", X"006C", X"0128", X"FFF2", X"FFA4", X"00CC", X"00AF", X"0193", X"00A5", X"FFBB", X"0355", X"04BA", X"052B", X"03EB", X"03ED", X"05BA", X"04D3", X"035C", X"0415", X"05E4", X"06A5", X"0715", X"03F5", X"05E3", X"0611", X"02DC", X"01D0", X"0346", X"013B", X"FFD4", X"0109", X"006E", X"FF66", X"00F9", X"0180", X"031A", X"0051", X"01EB", X"0247", X"01DA", X"036C", X"059F", X"0677", X"082A", X"07E1", X"0A77", X"0502", X"05E5", X"0832", X"0746", X"0503", X"058A", X"069F", X"0216", X"03ED", X"01E1", X"FF54", X"FFF0", X"0067", X"006E", X"000A", X"FF99", X"00AD", X"FE9C", X"FDB1", X"FCA1", X"FD48", X"FE07", X"FE73", X"FE6D", X"FCDE", X"FDB9", X"FAE2", X"0083", X"FF39", X"FF31", X"FD2C", X"FFC0", X"FF12", X"FFE6", X"FFD0", X"FFF2", X"FE7A", X"010E", X"003E", X"006A", X"006D"),
        (X"00FD", X"007D", X"FF69", X"FF3E", X"FFB6", X"FF04", X"FEC8", X"005A", X"0090", X"0066", X"003F", X"0054", X"0126", X"FF90", X"0036", X"00B7", X"0085", X"FFFE", X"0043", X"FFF8", X"FF4E", X"FFBC", X"FF05", X"0196", X"007B", X"FFE2", X"FF36", X"01A3", X"FFB3", X"FF68", X"FE8B", X"FF7C", X"010F", X"001F", X"FE92", X"FDD7", X"FF3A", X"FFBB", X"FE28", X"018D", X"011C", X"009A", X"FFFA", X"0376", X"0126", X"003E", X"000E", X"FEA8", X"FF4E", X"0185", X"FFEF", X"0030", X"0012", X"FF53", X"FFC8", X"FFFA", X"FF6F", X"001E", X"FFE9", X"03BA", X"014D", X"FFC9", X"002C", X"017F", X"FD31", X"FBD6", X"FBA5", X"FC0F", X"FEA9", X"FF0F", X"FDAF", X"FF47", X"01AE", X"00D7", X"0193", X"00E3", X"0060", X"0105", X"FFC6", X"019B", X"FEFB", X"FDE2", X"FFC4", X"FF7A", X"018C", X"FFBF", X"01BB", X"0070", X"FF80", X"FF00", X"FE67", X"FF29", X"FE13", X"FD74", X"FC76", X"FE8F", X"FEBB", X"FF91", X"011C", X"00A7", X"00BA", X"00EA", X"01AE", X"003B", X"015B", X"01A1", X"008C", X"0161", X"033F", X"01A6", X"00FC", X"FF1B", X"001E", X"FF03", X"0296", X"0314", X"FE8F", X"FDCD", X"FDA3", X"FFB5", X"FB8E", X"FB53", X"FA82", X"FE93", X"FE42", X"FF93", X"FF9D", X"0263", X"01A1", X"0338", X"0265", X"000F", X"FF64", X"FEE7", X"FEE8", X"FD53", X"00C9", X"02A2", X"0303", X"00F9", X"FFEE", X"FFF9", X"FF55", X"00CD", X"FCD5", X"FEF9", X"FD76", X"FE92", X"FC9D", X"FD8C", X"FE0C", X"013C", X"01FC", X"0567", X"0350", X"030C", X"039D", X"00F8", X"0372", X"00E3", X"0196", X"00AD", X"FE6F", X"FB5D", X"FDAA", X"0357", X"0185", X"FFF1", X"FFD1", X"0013", X"00A4", X"FF61", X"FBDA", X"FD77", X"FE6F", X"FDEE", X"0035", X"0057", X"01F2", X"04F4", X"082A", X"08AB", X"0A7B", X"077B", X"05AD", X"04A3", X"04AF", X"02EF", X"03CC", X"028F", X"0163", X"FE98", X"FE8F", X"FFC6", X"FE6C", X"0198", X"0058", X"002F", X"FE93", X"FFA3", X"FE7E", X"FE7C", X"00BA", X"FF8E", X"0256", X"0396", X"0416", X"037F", X"07C0", X"0815", X"0668", X"06CC", X"05CF", X"0413", X"040F", X"039D", X"0312", X"0387", X"00B0", X"02E5", X"FF69", X"FD31", X"FD24", X"038A", X"02C6", X"000A", X"008A", X"01BB", X"FED0", X"FEE3", X"00D1", X"0343", X"0465", X"0336", X"01DB", X"0319", X"056E", X"064C", X"07CE", X"0509", X"056B", X"01AB", X"02E5", X"00F1", X"00F8", X"01C7", X"01BB", X"009F", X"02EC", X"FE13", X"01B7", X"02BF", X"FFED", X"038F", X"0088", X"02D1", X"023E", X"FF42", X"0437", X"0426", X"030F", X"00BC", X"0104", X"0365", X"02E4", X"06B5", X"07B2", X"038B", X"00A4", X"FFE7", X"01FC", X"0103", X"FFDD", X"FDE0", X"005E", X"02F7", X"00A3", X"FF16", X"03A0", X"FE7E", X"024E", X"0009", X"03A2", X"014E", X"03D8", X"02B5", X"0500", X"043D", X"02E3", X"01C0", X"02B0", X"0403", X"0446", X"065C", X"0548", X"FF1F", X"FD0E", X"FE3E", X"FFB7", X"0178", X"00CD", X"0014", X"FFE4", X"0249", X"00B6", X"FEBC", X"00EF", X"031B", X"0030", X"0143", X"01E0", X"0159", X"046C", X"0448", X"04AC", X"045C", X"039B", X"052D", X"074D", X"0707", X"04ED", X"068E", X"03DF", X"000F", X"FD85", X"0273", X"03D4", X"0147", X"00D4", X"0183", X"044E", X"04FC", X"0316", X"03D3", X"056F", X"0323", X"0082", X"00F4", X"02E1", X"024A", X"05B9", X"05F0", X"062E", X"04F1", X"0194", X"03EC", X"032F", X"01DB", X"00C9", X"0181", X"05A3", X"0026", X"004B", X"03A2", X"01D4", X"00AD", X"02FC", X"0385", X"0538", X"0753", X"0278", X"0209", X"0261", X"0101", X"007C", X"02E0", X"025E", X"0433", X"05E7", X"02D9", X"03A6", X"0245", X"0152", X"0060", X"FD74", X"FA64", X"FA3B", X"FE77", X"002F", X"0096", X"FEAC", X"00B3", X"023C", X"01D0", X"014E", X"FF9E", X"0107", X"FF39", X"FDD8", X"FD7B", X"003F", X"FEE8", X"FEA1", X"004E", X"0257", X"FD0F", X"FF94", X"0060", X"FE55", X"FCAD", X"FC78", X"FBF5", X"FA74", X"F735", X"F6E3", X"FBE3", X"FE6D", X"FE53", X"FC9B", X"FE60", X"FEF8", X"FE05", X"FF24", X"010B", X"FEA4", X"FBC0", X"FBD6", X"FC8C", X"FC45", X"FEEB", X"FF52", X"00CF", X"FC25", X"F96B", X"FA39", X"FA81", X"FB36", X"FBB5", X"FBD3", X"FBE5", X"FB0F", X"F842", X"F922", X"FAD4", X"FC15", X"FCC5", X"FB96", X"FD17", X"FED3", X"FD0E", X"FF8F", X"FF24", X"FE1E", X"FEF1", X"FC18", X"FBC0", X"FB46", X"FE06", X"FE0A", X"002B", X"0195", X"FA9C", X"FAA5", X"F907", X"F950", X"FB4E", X"FBA4", X"FE2A", X"FD71", X"FC96", X"FB2C", X"FB7E", X"FCEA", X"FBB5", X"FB43", X"FC09", X"FB20", X"FC59", X"FCF4", X"FA8E", X"FD29", X"FE80", X"FA7E", X"F678", X"F8E4", X"FE74", X"FF2B", X"007C", X"FE69", X"FBD8", X"F9F1", X"F9C6", X"FA57", X"FBE4", X"FE27", X"FEE5", X"FC45", X"FE04", X"FF2E", X"FE93", X"FBD8", X"FCF1", X"FB7D", X"FC9A", X"FC96", X"FF6F", X"FE19", X"FC8C", X"FDB2", X"FD9E", X"FBD8", X"F8CD", X"FE48", X"FFE8", X"0116", X"FFF1", X"0053", X"FBBE", X"FA87", X"FC15", X"FD91", X"FB59", X"FEDE", X"FEF8", X"FFF6", X"FE48", X"FE28", X"FCE3", X"FB61", X"FC76", X"FAC7", X"FD53", X"FD91", X"022D", X"FEC3", X"FE9B", X"0080", X"FC5E", X"F9B4", X"F933", X"FCB2", X"FDB9", X"FF50", X"01F9", X"0418", X"FE98", X"FD24", X"FDDD", X"FE75", X"FF57", X"FDC8", X"FF06", X"FEE4", X"FE56", X"FFDB", X"FD0C", X"FBD7", X"FBCD", X"FAF9", X"FC58", X"FE99", X"020D", X"0098", X"00C0", X"024A", X"000A", X"FDA5", X"FA61", X"FBA9", X"FB69", X"FFAD", X"01CC", X"01B0", X"FE72", X"FD60", X"010C", X"017A", X"FF31", X"FC61", X"FD1E", X"FE63", X"FF79", X"FF64", X"FF9F", X"FE71", X"FE73", X"FD93", X"FEEC", X"FDE3", X"0139", X"00B4", X"021A", X"0474", X"0224", X"FFDF", X"FF40", X"FBC8", X"00A0", X"FE3E", X"0120", X"FFA0", X"FEA5", X"011C", X"017E", X"03AD", X"0154", X"00D2", X"0132", X"028B", X"03AC", X"0244", X"020D", X"0159", X"00C6", X"01EB", X"0085", X"FEBF", X"0159", X"021B", X"0186", X"01C2", X"0025", X"FFC0", X"FEAC", X"FAF4", X"0051", X"0032", X"0177", X"FF1F", X"FC85", X"FF52", X"000D", X"051F", X"040C", X"0216", X"04E8", X"0403", X"06B0", X"04FD", X"03BF", X"0526", X"0338", X"046A", X"0357", X"0383", X"00CF", X"0024", X"FFDB", X"035B", X"0268", X"022F", X"00A2", X"FD97", X"0082", X"FF53", X"FF53", X"FD5D", X"FFC9", X"00E1", X"FF0C", X"00A2", X"021E", X"046F", X"0333", X"04FE", X"03C0", X"00DA", X"01F9", X"036A", X"02F7", X"0400", X"0627", X"0365", X"0253", X"02A3", X"FFEF", X"037C", X"0364", X"03E6", X"FF77", X"FD3F", X"FFA0", X"00B9", X"FFB5", X"FF74", X"02D8", X"02A1", X"02B7", X"041F", X"0220", X"0480", X"044F", X"0637", X"0316", X"0370", X"FEEC", X"001E", X"01C8", X"0213", X"01EB", X"0195", X"012A", X"02A4", X"0239", X"0533", X"0493", X"00C1", X"FDFE", X"FD09", X"0043", X"0206", X"00C2", X"00CA", X"0334", X"04AF", X"071E", X"0751", X"06C6", X"06F7", X"0B3B", X"08A6", X"056B", X"0420", X"042E", X"0340", X"02D8", X"02D0", X"04A0", X"05E0", X"0635", X"037D", X"051D", X"0631", X"0211", X"00A5", X"FD6B", X"FDE0", X"FFFF", X"FF86", X"FFEB", X"FFD5", X"0120", X"03F7", X"05CC", X"0656", X"0951", X"0845", X"0833", X"0873", X"0925", X"0A54", X"0C8B", X"0F84", X"0A14", X"09AD", X"09BE", X"0C7A", X"09BB", X"0AC6", X"0726", X"04E1", X"01DD", X"02E1", X"000F", X"FF31", X"006F", X"0035", X"012E", X"001C", X"013A", X"FFDF", X"FFA4", X"03EC", X"0320", X"030E", X"04B6", X"04C0", X"0453", X"062E", X"0775", X"0964", X"05C6", X"0460", X"04EC", X"0623", X"054C", X"0368", X"0446", X"0339", X"FFCB", X"003E", X"FF01", X"006C", X"FF34"),
        (X"FEE2", X"004D", X"0006", X"000A", X"0076", X"009B", X"005C", X"012A", X"00F0", X"FFF4", X"FFCD", X"0162", X"FF7E", X"00C0", X"FEDE", X"0010", X"FE9F", X"00B6", X"001A", X"002F", X"FFDB", X"0018", X"01AB", X"FF2B", X"FEE8", X"FF7B", X"016B", X"0074", X"0021", X"010B", X"FFEF", X"0039", X"0080", X"FFCC", X"0171", X"0234", X"033B", X"03C9", X"01FC", X"0230", X"040D", X"03AA", X"035F", X"03F2", X"0026", X"0266", X"018F", X"01BE", X"014F", X"0069", X"017D", X"01D1", X"FF7C", X"FFA3", X"011D", X"FE86", X"0185", X"FECF", X"017B", X"01AB", X"0089", X"0134", X"03A8", X"042F", X"05AF", X"075E", X"07E5", X"0A17", X"0A8B", X"0A0E", X"0990", X"0607", X"006C", X"00D4", X"00E1", X"0042", X"FFFF", X"0095", X"024C", X"FFDE", X"014B", X"0056", X"0054", X"002A", X"FF8A", X"FFFE", X"00E6", X"FED7", X"000E", X"FF5D", X"009D", X"0182", X"02ED", X"03BC", X"0074", X"0220", X"013D", X"0391", X"FF7E", X"FF42", X"FF9E", X"FF22", X"FE32", X"0001", X"FF62", X"FE49", X"FFEB", X"024E", X"0049", X"02C3", X"00CC", X"0051", X"00C7", X"FFB4", X"FE39", X"FE16", X"FF2E", X"FE7E", X"FD4D", X"FEB4", X"0044", X"004D", X"FF5A", X"FE6E", X"0077", X"007E", X"FFFA", X"FDBA", X"FCC5", X"FC58", X"F9CC", X"FD8D", X"FF80", X"FCAE", X"FD64", X"012C", X"FCAB", X"FAF5", X"0172", X"027C", X"01DD", X"0127", X"008E", X"FE35", X"FF75", X"FB0A", X"FAE6", X"FC68", X"FF81", X"FD76", X"FB05", X"FCED", X"018B", X"0396", X"0467", X"00F8", X"FEBA", X"FF75", X"FEC4", X"0114", X"FFD3", X"0083", X"FF18", X"006B", X"FE3A", X"FC0E", X"FC84", X"0084", X"FF03", X"FF88", X"FEEA", X"FC46", X"00E3", X"F892", X"FCAB", X"FDB4", X"FC54", X"F90B", X"FA43", X"FC7B", X"FE68", X"FFFB", X"0277", X"0243", X"FFD4", X"FF8F", X"FED0", X"00AD", X"0092", X"FF8B", X"00B0", X"FF80", X"FCA0", X"FA72", X"FAA7", X"FFA1", X"0187", X"FD3F", X"004B", X"FA92", X"009E", X"FCF5", X"FC92", X"FCB1", X"FB1A", X"FD07", X"FCA6", X"FD11", X"FC54", X"FDB5", X"FE57", X"FFE2", X"003F", X"FD39", X"FEC4", X"FF71", X"FE6A", X"FF2A", X"FF35", X"0030", X"FD2B", X"FB3C", X"FCC8", X"FEC5", X"0220", X"FE52", X"FD7E", X"FBC5", X"0099", X"FF84", X"FFBF", X"FE7E", X"FD83", X"FDC2", X"FC1B", X"FCCD", X"010D", X"FF61", X"FEB8", X"00E2", X"FF98", X"00A3", X"0112", X"0113", X"FF24", X"FE8B", X"FE0D", X"FE3C", X"F910", X"F82D", X"FE69", X"0116", X"003B", X"FCDC", X"FF4D", X"FED1", X"01BA", X"FFBF", X"0085", X"FF1C", X"FE3B", X"0043", X"00AC", X"FDBF", X"FF25", X"FFB1", X"00C4", X"FE6E", X"018F", X"00AD", X"008E", X"0142", X"FEE1", X"FF5A", X"FCDA", X"FF4D", X"F935", X"F5D6", X"FC32", X"FC2A", X"FFBD", X"FD81", X"FF96", X"FB4E", X"00B9", X"0204", X"0032", X"FDF9", X"FE80", X"FE3C", X"FFDF", X"FE62", X"FE7D", X"FEBC", X"014F", X"FD53", X"FF02", X"00F6", X"0310", X"0351", X"01F0", X"00D8", X"0101", X"0338", X"FC8B", X"F5E9", X"F7CF", X"FCED", X"FF22", X"FEE0", X"FB25", X"FA78", X"FDE5", X"00CC", X"FEAF", X"FD1F", X"FC69", X"FFA9", X"FF4A", X"FE0C", X"FE0C", X"0037", X"00AD", X"FC9C", X"FD41", X"FE3D", X"0078", X"0362", X"0403", X"05FA", X"06FE", X"0924", X"0799", X"FBE5", X"F955", X"FED4", X"FF96", X"FDBC", X"FB0A", X"FCA9", X"FDE5", X"FE11", X"008F", X"FCED", X"FD71", X"FDFF", X"FD57", X"FDCF", X"0111", X"0182", X"01E6", X"FE56", X"FD10", X"FE78", X"FE7F", X"00B8", X"FF61", X"0326", X"0579", X"0887", X"0C38", X"0465", X"FB22", X"00F6", X"0151", X"FDE8", X"FC48", X"FDFD", X"FCAB", X"FED7", X"0042", X"FD46", X"FC47", X"FBC8", X"FCE5", X"FE1C", X"FF71", X"FEB6", X"001B", X"00D1", X"FDDE", X"FD32", X"FE54", X"FF3E", X"FDFD", X"FEA7", X"003F", X"0554", X"0795", X"0477", X"01AA", X"02B0", X"FE50", X"FD8D", X"FC91", X"FD5E", X"FEDF", X"036F", X"0419", X"01CD", X"0063", X"FDD4", X"FDE9", X"FE56", X"FB5C", X"FDD8", X"FFC9", X"0003", X"FD33", X"FEA4", X"FEA5", X"FF35", X"FDDD", X"FCFA", X"FD8D", X"FDA7", X"00AB", X"076B", X"0292", X"034A", X"008E", X"FE92", X"FDB9", X"FBDA", X"03E8", X"0775", X"084E", X"0832", X"05AF", X"0277", X"0128", X"FE22", X"F99D", X"FE28", X"00D5", X"FF08", X"FDFD", X"FF18", X"FF26", X"0051", X"004C", X"FE12", X"FD21", X"FBB3", X"FD15", X"068F", X"0236", X"027F", X"00BC", X"FE8E", X"FDC4", X"FE32", X"058A", X"0A05", X"0CA8", X"0E0D", X"0E58", X"0A79", X"0842", X"0677", X"00CC", X"003E", X"015A", X"FFFB", X"FFC1", X"0059", X"FF8A", X"0014", X"00C1", X"FF88", X"FD49", X"FE6D", X"FD7B", X"0727", X"04DE", X"040A", X"FFBA", X"FE3A", X"FECB", X"FC99", X"020D", X"069B", X"0A37", X"0B2C", X"0D6C", X"10A7", X"101C", X"0DBF", X"0BFB", X"0763", X"0510", X"FF85", X"FF53", X"FE20", X"FFD1", X"000F", X"038D", X"0114", X"015D", X"FE5B", X"FD35", X"06E6", X"02CB", X"011F", X"FEAD", X"FE96", X"FDFC", X"F88F", X"006F", X"00E3", X"02BB", X"04E0", X"066E", X"08BD", X"0BDC", X"0DF9", X"0C2A", X"07BC", X"0281", X"FF29", X"FE64", X"FDE0", X"01D1", X"FFEC", X"00BA", X"0082", X"0293", X"0135", X"0095", X"04CD", X"FE21", X"0080", X"0100", X"FDEA", X"FD8C", X"F79E", X"FC80", X"FE92", X"FDC8", X"FE36", X"FED1", X"00C3", X"01CA", X"03E5", X"0785", X"055E", X"012D", X"0169", X"0186", X"0078", X"0156", X"0059", X"0198", X"02CC", X"0369", X"01E8", X"FEC6", X"0296", X"02B9", X"0111", X"FED9", X"FF16", X"FE0B", X"F98F", X"FC86", X"FCB5", X"FE93", X"FDBE", X"FDC3", X"FD15", X"FF15", X"FF70", X"01D9", X"01E9", X"0191", X"0262", X"0103", X"0040", X"FF73", X"01B4", X"0086", X"0163", X"0081", X"0138", X"FF25", X"012D", X"029F", X"FF75", X"0156", X"FE46", X"FDA5", X"FD10", X"FCC9", X"FDC4", X"FF24", X"FEE1", X"FD44", X"FE94", X"FEBA", X"FF82", X"FF1F", X"00FD", X"0113", X"0331", X"0051", X"FF6A", X"00E8", X"FFDC", X"0066", X"FFB1", X"0173", X"0343", X"0006", X"01EB", X"0201", X"FEE9", X"FF3E", X"007C", X"FED5", X"FC18", X"FE25", X"01E5", X"02B8", X"0152", X"007E", X"FFF9", X"FFA3", X"003E", X"0054", X"0000", X"00F9", X"014C", X"0044", X"00D2", X"0074", X"FF48", X"00F9", X"025A", X"0309", X"032F", X"0313", X"0144", X"012F", X"0016", X"0066", X"FE67", X"FC73", X"F9ED", X"F81A", X"FC73", X"FF9F", X"FFD6", X"0086", X"00C1", X"FE88", X"0144", X"038C", X"02B8", X"035D", X"04A7", X"03A1", X"011F", X"0154", X"019B", X"0069", X"FF96", X"04B9", X"0411", X"FF98", X"02B4", X"FE09", X"FFE1", X"FF35", X"00CE", X"FEC7", X"F79B", X"F54F", X"F5D9", X"F880", X"F8D4", X"FE44", X"FCE6", X"FDD8", X"FEBB", X"02AE", X"02B4", X"026F", X"02C1", X"0216", X"FEA0", X"FEBA", X"FE25", X"FB29", X"FC4F", X"FD41", X"FF80", X"FFA5", X"03E3", X"0101", X"FEA4", X"0081", X"0150", X"FF77", X"FDF3", X"F8DA", X"F244", X"F442", X"F47F", X"F40D", X"F374", X"F386", X"F657", X"F53B", X"F708", X"F5BF", X"F699", X"F4FA", X"F415", X"F5F4", X"F727", X"F629", X"F4E3", X"F7E3", X"F9C8", X"FB43", X"00B3", X"01AB", X"00C7", X"FF0A", X"00F5", X"FF7B", X"000A", X"FCF5", X"F96C", X"F9ED", X"FCE9", X"FBF3", X"F72D", X"F78A", X"F96C", X"FABF", X"F75E", X"F765", X"F5C3", X"F5E9", X"F622", X"F902", X"FB11", X"F9E7", X"FA0B", X"FB12", X"FBDA", X"002C", X"FF94", X"00A4", X"FFB3", X"FFF1", X"0008", X"0054", X"FFF8", X"FE61", X"FE4A", X"FFA3", X"0108", X"FF56", X"FF16", X"FDE1", X"FD34", X"FE0A", X"FC52", X"FD54", X"FC46", X"FCBE", X"FD19", X"01F8", X"FFB9", X"FE68", X"FD74", X"FCF9", X"FD44", X"FF58", X"009F", X"017E", X"FF40"),
        (X"FFDB", X"FF76", X"009C", X"00B6", X"002D", X"FF9F", X"FEB5", X"FFC6", X"FFCB", X"0065", X"006C", X"0073", X"FE79", X"FF79", X"0204", X"0005", X"00A1", X"FFCE", X"FF62", X"0076", X"FEF9", X"01EA", X"FEC0", X"0097", X"0086", X"FFE6", X"FEEE", X"FFA9", X"00F8", X"FF95", X"FEDF", X"FFE9", X"FF06", X"FFE2", X"FD81", X"FBE4", X"FD99", X"FE94", X"FD9B", X"FCAE", X"FB77", X"FD92", X"001F", X"0141", X"04DA", X"01D6", X"FE6A", X"FD55", X"FD32", X"FE7E", X"FEE1", X"FF2A", X"FE98", X"0074", X"FFCC", X"FFB8", X"015D", X"FFF8", X"0102", X"FFD2", X"FE95", X"FD57", X"FD19", X"FCC3", X"FC20", X"00C5", X"FFAF", X"0176", X"03D9", X"0165", X"FFD1", X"01D3", X"0555", X"033C", X"01E8", X"FF0E", X"FF1A", X"FBD0", X"FA8D", X"FECE", X"03FC", X"024D", X"FF64", X"FFEF", X"003D", X"00A8", X"0329", X"FFD7", X"FFB7", X"0247", X"02E1", X"0378", X"025F", X"0343", X"0356", X"0621", X"093F", X"0604", X"04AF", X"0315", X"02C2", X"00FE", X"00A4", X"005D", X"FFF3", X"FD73", X"F98E", X"F76C", X"FC45", X"FEDB", X"FD5A", X"FEC3", X"FF1B", X"FE03", X"0136", X"00B8", X"01F6", X"0508", X"07CB", X"035B", X"0286", X"02AC", X"069A", X"04A0", X"03A6", X"04AF", X"0295", X"0263", X"0273", X"FF69", X"0228", X"0187", X"FF6B", X"FE21", X"FD49", X"FD60", X"FC89", X"FFC4", X"FF5C", X"FE70", X"001E", X"FDCA", X"03A3", X"0517", X"0700", X"0888", X"0549", X"0241", X"0455", X"0248", X"0166", X"FF49", X"FF0F", X"FFD4", X"FF19", X"01DA", X"00A4", X"FE60", X"0168", X"0143", X"006F", X"003C", X"023D", X"0034", X"00B2", X"FF4A", X"016A", X"FC88", X"003C", X"0237", X"FF3B", X"042A", X"0627", X"0422", X"0210", X"010F", X"000E", X"0153", X"01F5", X"008E", X"00CF", X"0173", X"0275", X"FFBE", X"010A", X"0143", X"026E", X"FF55", X"02CF", X"01B7", X"0094", X"003E", X"020B", X"0286", X"0692", X"0011", X"FF06", X"01B6", X"FEA7", X"0164", X"04EB", X"0240", X"013C", X"012E", X"FFFA", X"0262", X"001D", X"0150", X"0301", X"044F", X"0487", X"00CA", X"018D", X"033F", X"02CD", X"02B9", X"018E", X"0145", X"018F", X"FDDF", X"FEB8", X"0425", X"0732", X"01E2", X"FE84", X"00BA", X"FF70", X"0152", X"01ED", X"008F", X"FF51", X"025C", X"015F", X"002E", X"028B", X"0286", X"0304", X"019F", X"0288", X"020A", X"00D5", X"0122", X"01D5", X"FFB3", X"FF9F", X"012C", X"006A", X"FF1B", X"001F", X"0719", X"0803", X"0353", X"00EC", X"FFEE", X"01FA", X"00E0", X"053F", X"014C", X"02D9", X"03E1", X"02A8", X"027A", X"FF85", X"FEDB", X"FEE0", X"FD7E", X"002F", X"00FF", X"008F", X"FD6A", X"FD0F", X"FB37", X"FDB3", X"FF77", X"FEB8", X"FE54", X"FF12", X"05C3", X"02B8", X"02C3", X"00F1", X"0065", X"025B", X"054B", X"0276", X"0384", X"0177", X"FEA0", X"FF35", X"FC9B", X"FB08", X"FABB", X"F96E", X"FACB", X"FDE3", X"FE5D", X"FD1C", X"FD0E", X"FBEC", X"FC1D", X"FB2A", X"FA74", X"FA61", X"F908", X"FA5F", X"040C", X"0245", X"0238", X"FFDC", X"FF72", X"0225", X"0085", X"0176", X"FDDA", X"FA25", X"F6CD", X"F757", X"F8E4", X"F948", X"FB53", X"F7C8", X"F96C", X"FBB1", X"FDDA", X"FE08", X"FCC5", X"FC7D", X"FDE7", X"FCFC", X"F659", X"F4D9", X"F28A", X"F3F1", X"FF40", X"FFD3", X"0176", X"FFF0", X"FCFF", X"FF80", X"FDB5", X"FE7D", X"F78B", X"F258", X"F296", X"F6FD", X"F8E9", X"FD2C", X"FC13", X"FC36", X"FB7C", X"FCEF", X"FE32", X"FC97", X"FC15", X"FE6B", X"FE21", X"FA44", X"F6F9", X"F481", X"EF84", X"F2A3", X"FE39", X"01F0", X"0266", X"FFED", X"FD33", X"FD9E", X"FCF7", X"F9DB", X"F440", X"F1B7", X"F534", X"F91F", X"FC24", X"0030", X"FE2C", X"FCE7", X"005C", X"0374", X"FE25", X"FCC5", X"FD98", X"0096", X"02A7", X"FCD2", X"F9B4", X"F641", X"F451", X"F73A", X"010F", X"04AB", X"00BC", X"014C", X"FF4D", X"FF8F", X"FE95", X"FB8D", X"F6FB", X"F886", X"F972", X"FD9C", X"00BA", X"FE25", X"FB10", X"FFAB", X"0317", X"02E3", X"0097", X"FCC8", X"FC0B", X"0088", X"FEA2", X"FE9B", X"FCE5", X"F9EC", X"FBB0", X"FE14", X"0488", X"078F", X"02D4", X"FF04", X"00B2", X"02D2", X"0225", X"0014", X"FE0E", X"FCB9", X"FDA9", X"FDCA", X"FF92", X"FDC3", X"FE49", X"0028", X"0360", X"0221", X"FFF3", X"FC3B", X"FB94", X"FDBD", X"003D", X"004F", X"FFA9", X"FE1C", X"FF92", X"051E", X"08E5", X"0811", X"0343", X"FEE0", X"00FF", X"03E8", X"06B5", X"04AA", X"0157", X"FDF4", X"FA2A", X"F70C", X"FA3A", X"FD1E", X"FC0F", X"FE0D", X"02FA", X"0178", X"FD40", X"FACA", X"FDE8", X"FFDD", X"025B", X"0172", X"027A", X"02C0", X"04C0", X"081B", X"0C6D", X"0981", X"03CA", X"FF15", X"01F9", X"036A", X"0A57", X"065E", X"03FE", X"0033", X"FA30", X"F6E8", X"F67B", X"F718", X"F640", X"F8CD", X"FF65", X"00B7", X"FC48", X"FD12", X"FEA8", X"0063", X"01D0", X"02DA", X"04AB", X"03D5", X"05B0", X"06B2", X"0BD0", X"08AF", X"03A0", X"FEF9", X"00A4", X"00B6", X"0A1A", X"08D2", X"05C8", X"00FA", X"FB8D", X"FB9A", X"F8CE", X"F7AB", X"F513", X"FA5B", X"FF15", X"0016", X"0075", X"01AC", X"0348", X"04D2", X"03F7", X"0022", X"0431", X"032E", X"0395", X"07DD", X"0A93", X"05C4", X"0360", X"0119", X"0035", X"01F8", X"0788", X"067A", X"067C", X"02AF", X"0272", X"FFEB", X"FDBA", X"FDA2", X"FC5A", X"FC60", X"0330", X"020C", X"02E6", X"0430", X"0420", X"038D", X"0236", X"0310", X"0375", X"0242", X"0262", X"03D8", X"080B", X"06BB", X"0235", X"00B9", X"00F5", X"00EA", X"07CE", X"0642", X"03D2", X"05FF", X"035B", X"04CC", X"0558", X"0397", X"05AF", X"006F", X"FEC9", X"01B7", X"0337", X"04BE", X"0451", X"0587", X"024E", X"02AD", X"027B", X"0096", X"014F", X"03CD", X"08C9", X"055F", X"01CB", X"016E", X"01E8", X"04C4", X"07C6", X"06B3", X"031D", X"04AF", X"04AA", X"0475", X"0403", X"0418", X"0267", X"00DB", X"FE66", X"0150", X"02D7", X"03F1", X"023A", X"04BD", X"0427", X"01DD", X"02E3", X"FF85", X"02B1", X"0660", X"06D9", X"0597", X"01AA", X"00CB", X"0110", X"05C0", X"0712", X"063C", X"04A8", X"01FD", X"024B", X"021D", X"03CC", X"02A6", X"0124", X"FD66", X"FE2E", X"FF63", X"0013", X"01C0", X"0297", X"058D", X"06A0", X"03F5", X"030D", X"0369", X"0498", X"0605", X"0458", X"FF42", X"005A", X"FFB6", X"FF5B", X"0299", X"05B7", X"07FE", X"05E4", X"03C3", X"02C8", X"FFEA", X"00FD", X"01E2", X"012D", X"FE20", X"FDE0", X"FDA4", X"FE2D", X"FF5F", X"0449", X"02C2", X"034E", X"006C", X"02C7", X"0416", X"044E", X"02FF", X"04CC", X"03AA", X"00E1", X"FFA1", X"0124", X"0056", X"03DF", X"07A1", X"01D5", X"04A7", X"01FF", X"0036", X"00FC", X"0276", X"02CF", X"0034", X"013F", X"01DD", X"FF18", X"001C", X"02DA", X"014F", X"FFA6", X"FE8C", X"00F4", X"028D", X"015C", X"050D", X"05C8", X"0449", X"FF67", X"0166", X"FF3A", X"010B", X"FE11", X"0092", X"00C7", X"0045", X"010E", X"037D", X"031F", X"0399", X"0225", X"04BC", X"0296", X"FF82", X"FC83", X"FCA2", X"FE1E", X"FCDB", X"00A7", X"FC8A", X"FC65", X"FDD0", X"FFEC", X"028D", X"02AB", X"01C0", X"014C", X"002D", X"FF5D", X"FEBE", X"FE92", X"FD4D", X"FE83", X"FCC3", X"FB8E", X"FBB2", X"F83F", X"FAEC", X"FC38", X"FC42", X"FCC4", X"FB22", X"FDBC", X"FF87", X"FE84", X"00CD", X"0063", X"FE8F", X"FD2F", X"FCD1", X"FF0B", X"009B", X"0115", X"FFC7", X"015F", X"0153", X"007B", X"0076", X"000D", X"00E1", X"FF83", X"018D", X"0009", X"0015", X"01BD", X"FE6F", X"0126", X"0003", X"005C", X"FD62", X"FE3D", X"FE75", X"FCBA", X"FCF9", X"FC7A", X"FECE", X"FE2C", X"FD50", X"008B", X"FED8", X"FDC6", X"FF1A", X"FFA9"),
        (X"003F", X"FEF7", X"FF49", X"FF3D", X"FFD4", X"00BF", X"FF4A", X"FFA4", X"0142", X"001C", X"000B", X"0053", X"FDC7", X"FE22", X"FFBD", X"00DA", X"0044", X"FFD4", X"FFD3", X"006B", X"0021", X"FF8F", X"00AD", X"FEFA", X"017F", X"007B", X"001B", X"FFC1", X"016A", X"FFD0", X"FDFD", X"0041", X"FF86", X"FF9E", X"FD62", X"FCFF", X"FD4B", X"FB49", X"FC1E", X"FFE3", X"FF64", X"FEB8", X"FFC6", X"FA92", X"FCAA", X"FE0E", X"FA32", X"FD1A", X"F8D5", X"FB08", X"FC48", X"FD4D", X"FFA4", X"01A2", X"FFD6", X"013C", X"00F4", X"0147", X"FF77", X"FF8B", X"FDB6", X"FE2A", X"FC35", X"FA99", X"F8BC", X"F739", X"F4AB", X"F672", X"F57D", X"F9F9", X"FAD8", X"F75C", X"F704", X"F6F2", X"F736", X"F609", X"F529", X"F340", X"F6EB", X"F88D", X"FBDB", X"FDAA", X"FFA2", X"FF7F", X"0016", X"006A", X"FF4A", X"FF2A", X"0048", X"FC60", X"F9CA", X"F6B4", X"F6B1", X"F4A3", X"F710", X"F631", X"F5DF", X"F54B", X"F7C9", X"F69A", X"F53C", X"F349", X"F1E4", X"F6C1", X"F811", X"FAE5", X"023A", X"0167", X"029C", X"FE7A", X"FF86", X"FF7E", X"FEF7", X"0082", X"FD6D", X"FC5B", X"FC42", X"FB09", X"FA34", X"FB03", X"F9D2", X"FA5C", X"FB0C", X"FD7C", X"FEB5", X"FD71", X"FEC6", X"0087", X"0095", X"01DF", X"FF23", X"00D3", X"0230", X"075D", X"0678", X"09AF", X"0623", X"0226", X"FE54", X"FFD3", X"FF90", X"0096", X"FE37", X"FEE8", X"FADB", X"FB57", X"FB69", X"FD0F", X"FB81", X"FDE8", X"FC66", X"FDBC", X"FC72", X"FCB1", X"FF63", X"0142", X"04E0", X"0621", X"052F", X"063A", X"07BA", X"0AEB", X"0C09", X"0D9E", X"09E0", X"0633", X"0334", X"0127", X"0015", X"006A", X"FF82", X"FA8F", X"FC50", X"FF45", X"FEBC", X"FF96", X"FF25", X"FEB6", X"FD71", X"FD18", X"FC9E", X"FB23", X"FAD0", X"FD1E", X"FE0D", X"FDED", X"0113", X"04DF", X"0638", X"07A7", X"0C4A", X"0E97", X"0C23", X"0826", X"0312", X"003B", X"006B", X"FD14", X"FE52", X"FACC", X"FAD6", X"0201", X"01BE", X"00B6", X"01B0", X"FF44", X"FD11", X"FC9B", X"FBF3", X"FBA3", X"FA76", X"FB80", X"FD70", X"00E9", X"0281", X"0312", X"02BC", X"05A3", X"0AB2", X"0EA4", X"0E18", X"09E7", X"0486", X"0110", X"0179", X"FC8E", X"FF2B", X"FBFB", X"FB31", X"00F8", X"0216", X"019D", X"00FF", X"00AF", X"FF21", X"FD8A", X"FD78", X"FAB3", X"FAC9", X"FCC9", X"013C", X"0172", X"FFC4", X"00B6", X"01FB", X"031B", X"046D", X"0B88", X"0F51", X"097A", X"025F", X"004D", X"FF3F", X"FD7F", X"FE8B", X"FB6B", X"F9E9", X"FF9C", X"FEE8", X"0032", X"01B0", X"0179", X"FFB7", X"00A2", X"01C7", X"FDF1", X"F867", X"FCB0", X"009E", X"0199", X"01D4", X"014D", X"0031", X"025B", X"022C", X"040F", X"0C1F", X"078F", X"00AF", X"FEA2", X"FFFA", X"FD4C", X"FC5B", X"FB63", X"001B", X"FE92", X"FD24", X"FFE8", X"01A5", X"043E", X"037E", X"0570", X"0449", X"FE51", X"F8B5", X"FEA8", X"0243", X"00F6", X"FF8A", X"0000", X"0018", X"0081", X"FF2A", X"0109", X"063B", X"0962", X"0328", X"0150", X"0005", X"FD3C", X"F902", X"FB66", X"FC02", X"FE2C", X"003E", X"009F", X"0272", X"044B", X"04D8", X"04B9", X"0627", X"01F3", X"FA0D", X"FFDC", X"0171", X"FD86", X"FC60", X"FE1E", X"FA89", X"FC87", X"FD21", X"FD23", X"001D", X"0316", X"05FE", X"01A3", X"FFBC", X"FDAA", X"FAEC", X"FC24", X"FB19", X"0168", X"0317", X"02D4", X"0249", X"0332", X"05EE", X"0852", X"0ADA", X"02D4", X"FAE7", X"FD0B", X"FD9B", X"FB0F", X"FBA8", X"FEA6", X"FD1E", X"FE6E", X"FC3E", X"FB19", X"FDF5", X"FECF", X"FF62", X"FCBA", X"FEEC", X"00C3", X"FA23", X"FAEB", X"FEA3", X"03E1", X"042D", X"0159", X"0271", X"041F", X"055D", X"0952", X"090C", X"FF72", X"F9F1", X"FC3B", X"FC3F", X"FB99", X"FD03", X"0083", X"02EE", X"FE11", X"FEE1", X"FC98", X"FC83", X"FBDA", X"FB9C", X"FCCA", X"030C", X"FE19", X"FD88", X"FB36", X"02D2", X"0608", X"018C", X"042E", X"03B3", X"035F", X"0577", X"072A", X"02A1", X"FE59", X"FBB6", X"FC82", X"FBD9", X"FE6D", X"FF46", X"008C", X"00A6", X"FE4E", X"FD1C", X"FF2E", X"00D8", X"FD75", X"F7F3", X"FDEC", X"02A2", X"FDA9", X"0095", X"FBC2", X"05EF", X"043A", X"026D", X"0373", X"05A2", X"05C7", X"05E2", X"0272", X"0145", X"FE64", X"FEDF", X"FDCD", X"FEAB", X"FE2D", X"FEFA", X"FE66", X"FD7E", X"FE70", X"FC64", X"00C0", X"FE58", X"FA40", X"FBD2", X"FC83", X"FDA2", X"FDA3", X"FC7A", X"FB3A", X"0023", X"037A", X"0221", X"026A", X"0459", X"0504", X"0214", X"FEBA", X"FF96", X"FEEE", X"FFC2", X"0173", X"FF12", X"FFAE", X"FE1F", X"FE3D", X"FF45", X"FE5C", X"FE33", X"00CE", X"FF83", X"F7CF", X"FA94", X"FD95", X"0054", X"FF21", X"FC46", X"FB95", X"FFE9", X"04CA", X"0329", X"020F", X"023E", X"05E2", X"025D", X"FE6A", X"FF02", X"FFA2", X"013A", X"0189", X"0091", X"FF1D", X"FD4E", X"FE00", X"00E7", X"0003", X"FFFF", X"0098", X"00C9", X"F655", X"F8F7", X"FF90", X"FCBF", X"FDEB", X"FC64", X"FB5A", X"0116", X"0309", X"030E", X"0283", X"0417", X"0500", X"00A1", X"FF6A", X"FEBE", X"00AF", X"FFC6", X"FF32", X"FE29", X"FCD7", X"FC96", X"FF5F", X"FEFF", X"FF44", X"FE29", X"FE5C", X"00FF", X"F957", X"FA8F", X"FC0E", X"FED4", X"FFD4", X"00F6", X"FB8F", X"FEC5", X"0227", X"02FA", X"015C", X"0325", X"0261", X"FFCD", X"FD8E", X"FDC9", X"FCED", X"FE74", X"003E", X"FE24", X"FD60", X"FCCB", X"FE9B", X"FEE5", X"FF5A", X"FE5F", X"FF3E", X"FF62", X"FB4B", X"F99F", X"FBEF", X"001E", X"0221", X"FDF8", X"FAE6", X"FC1E", X"FD33", X"0192", X"FFFF", X"007C", X"FF89", X"00D2", X"FFB2", X"FD33", X"FCB9", X"FE0D", X"FEDF", X"FE61", X"00D0", X"FE3C", X"FCF0", X"FE00", X"0143", X"01A9", X"FEFB", X"FC0F", X"FBC2", X"FCDF", X"FEF4", X"FF0A", X"0008", X"FCD5", X"F99D", X"FC08", X"FE06", X"FFDB", X"0185", X"0071", X"0072", X"FF63", X"010D", X"0110", X"FD45", X"FE28", X"0119", X"009B", X"0036", X"012D", X"FE07", X"005F", X"036A", X"03F2", X"009F", X"FDFC", X"FF51", X"0321", X"002C", X"FEAB", X"004A", X"F928", X"FCB0", X"FCB5", X"FE1F", X"FFF1", X"00AC", X"FFEA", X"FE8F", X"00EA", X"0320", X"01EB", X"02CC", X"01E4", X"013C", X"02AF", X"01ED", X"01D7", X"017C", X"0191", X"0467", X"0289", X"0098", X"FF9F", X"0237", X"0271", X"FF91", X"FEEA", X"0099", X"FBCE", X"FE1B", X"FBA9", X"FDDB", X"FE9D", X"FFCC", X"005E", X"019C", X"0360", X"0575", X"04E6", X"0421", X"0497", X"03A8", X"02F2", X"01E0", X"01B6", X"00F0", X"0228", X"004F", X"007F", X"FFA9", X"FFD8", X"0476", X"0210", X"FF3B", X"FF31", X"FEC6", X"FF2B", X"FF7F", X"F9BE", X"FB21", X"FBC3", X"FD18", X"FFA2", X"006C", X"FEAF", X"0099", X"FE35", X"FE9F", X"FFAE", X"FD5F", X"FDC5", X"FE18", X"020B", X"01FB", X"005C", X"FED5", X"0120", X"FFD1", X"FCF9", X"FE49", X"FF16", X"0085", X"FFCE", X"0101", X"FE7A", X"02A2", X"FCCD", X"F5ED", X"F989", X"FA4C", X"F79E", X"FA69", X"F9AF", X"F956", X"F882", X"F9E7", X"FA7B", X"FC3B", X"FB6D", X"FB3A", X"FBF2", X"FA70", X"F783", X"FB45", X"FFBC", X"00E9", X"0035", X"002D", X"0071", X"FF19", X"FF84", X"FF8E", X"FE65", X"FF23", X"FA7C", X"F970", X"F69B", X"F51A", X"F330", X"F3EA", X"F415", X"F6F1", X"F716", X"F5C6", X"F216", X"F5D6", X"F674", X"F60B", X"F6AA", X"F6E7", X"F776", X"FB3F", X"FD9B", X"FEC6", X"FF90", X"FFBF", X"FF5C", X"FF94", X"00F4", X"00AA", X"FFFA", X"FF57", X"FF8C", X"002C", X"FC6A", X"FCCA", X"FB68", X"FA08", X"F7FF", X"FBAE", X"F79A", X"F97D", X"F7D7", X"F74D", X"F7C8", X"F8DE", X"F7E4", X"F98D", X"FC3A", X"FBDF", X"FA98", X"FE76", X"FF34", X"FF76", X"FF2A", X"004B"),
        (X"FEA2", X"0014", X"0201", X"0033", X"FFEB", X"FFEC", X"FF78", X"003C", X"FFFD", X"00A9", X"0139", X"FF5F", X"005E", X"0002", X"003D", X"002D", X"FF8E", X"FF87", X"0119", X"FF61", X"FFBC", X"0183", X"001A", X"FFAF", X"0096", X"FF77", X"0012", X"FF93", X"0014", X"FFCB", X"00B3", X"013F", X"01CB", X"0118", X"00F4", X"FFFF", X"02BB", X"0050", X"00AB", X"021A", X"007A", X"0102", X"FDB3", X"FE20", X"011D", X"0205", X"0139", X"FF12", X"0009", X"011C", X"FFF4", X"FF74", X"FF6B", X"0036", X"0027", X"FF57", X"000F", X"FE97", X"FFCD", X"FF31", X"FEA8", X"018D", X"000D", X"FFBF", X"038E", X"03D5", X"03E4", X"0429", X"04CE", X"0212", X"FF64", X"FF28", X"0166", X"052D", X"055C", X"04D1", X"030E", X"02FB", X"03BD", X"0201", X"0190", X"0312", X"0102", X"FF57", X"001F", X"FF32", X"FE79", X"FEA8", X"0052", X"02E1", X"0161", X"027C", X"05B9", X"01FC", X"05FA", X"0722", X"0889", X"0574", X"08B5", X"069D", X"073B", X"074F", X"0907", X"072D", X"0639", X"061A", X"056F", X"064F", X"052F", X"0273", X"03DC", X"FFC1", X"0155", X"FFA0", X"FD92", X"FE84", X"00EB", X"0278", X"0198", X"018E", X"04B4", X"0272", X"FFCD", X"0192", X"0232", X"013C", X"032A", X"0273", X"03E2", X"0555", X"0486", X"006B", X"00C1", X"00A1", X"007F", X"0045", X"0514", X"07C8", X"048F", X"0281", X"FF64", X"0015", X"FE78", X"FC64", X"FE41", X"0354", X"04BA", X"050D", X"0938", X"06C8", X"0405", X"0362", X"0267", X"02BB", X"0264", X"0224", X"040E", X"05EC", X"02A1", X"02D4", X"0224", X"FE89", X"FD3F", X"FED7", X"014B", X"0880", X"0333", X"026F", X"FF99", X"00C2", X"00E6", X"FDB0", X"FF18", X"0634", X"0741", X"0976", X"0A4F", X"0895", X"049C", X"01FD", X"02CB", X"0503", X"049D", X"05BB", X"04A6", X"040A", X"0190", X"0203", X"0048", X"FEED", X"FF46", X"FF1D", X"0259", X"0A52", X"042A", X"0048", X"0042", X"0248", X"0286", X"0242", X"02CD", X"04CD", X"082A", X"09C3", X"0A92", X"07B7", X"03F4", X"0179", X"03EA", X"0335", X"0253", X"042C", X"03D9", X"0245", X"00DC", X"FFDA", X"0049", X"00C6", X"FEFA", X"00E0", X"0777", X"091C", X"035A", X"03DA", X"0035", X"02F0", X"0128", X"00D7", X"0135", X"0341", X"070E", X"0879", X"080D", X"0705", X"0411", X"01B3", X"00A3", X"FFE4", X"FFEA", X"0024", X"0006", X"FEF0", X"01CE", X"01D0", X"0297", X"02B9", X"0257", X"052B", X"083E", X"08AE", X"04F7", X"023C", X"0103", X"000F", X"027F", X"021F", X"0525", X"0481", X"0618", X"04B4", X"07DB", X"0853", X"044F", X"01A1", X"FF7A", X"FE8F", X"FE0D", X"FC4D", X"FE3D", X"FFAF", X"01DC", X"040C", X"05F8", X"029A", X"04E2", X"07C5", X"08B1", X"071A", X"033B", X"02FE", X"FFBE", X"FEF8", X"00AE", X"0397", X"036A", X"0589", X"0791", X"0804", X"0775", X"0703", X"021A", X"FF0A", X"FF39", X"FCB6", X"FB7F", X"F714", X"FB81", X"004C", X"029E", X"02DC", X"05BF", X"0587", X"0939", X"07E6", X"0923", X"03B5", X"0330", X"FE75", X"FFD7", X"001F", X"0024", X"0404", X"015B", X"00A5", X"05B0", X"0725", X"08A7", X"05BB", X"039D", X"FF95", X"FD7B", X"FC02", X"F9B0", X"F95A", X"FB97", X"FFDD", X"0013", X"0231", X"057B", X"0844", X"08F4", X"08C1", X"0880", X"0411", X"0179", X"FF4B", X"FFF6", X"014B", X"032D", X"FFB9", X"FE87", X"0463", X"03E8", X"0780", X"0690", X"050A", X"0339", X"FF70", X"FC66", X"FAD5", X"F9E7", X"FAB2", X"FC68", X"FF4A", X"0330", X"04C4", X"04F4", X"0527", X"0383", X"03D5", X"05BC", X"064C", X"080D", X"00F3", X"000B", X"00D0", X"021F", X"FD6A", X"FF90", X"036C", X"02C7", X"0334", X"03F5", X"0354", X"01B6", X"FF1E", X"FD47", X"F9C2", X"FB1E", X"FBC1", X"FC83", X"FDE7", X"0277", X"0652", X"0636", X"0381", X"04E6", X"0568", X"06CE", X"062C", X"0499", X"01D2", X"FF2B", X"01E8", X"FDAC", X"FD0A", X"FD59", X"051E", X"038D", X"0295", X"025B", X"03E6", X"0243", X"FF94", X"FE29", X"FAB7", X"FB28", X"FBBE", X"FC96", X"03BD", X"079B", X"0803", X"07CD", X"030A", X"0304", X"0213", X"0239", X"043F", X"0500", X"0060", X"008E", X"004B", X"FE26", X"FF37", X"002B", X"0660", X"0673", X"03B6", X"01C9", X"0196", X"FF87", X"FE99", X"FCFD", X"FAB6", X"FC23", X"FD33", X"FECD", X"0722", X"075F", X"0806", X"0773", X"040F", X"0486", X"0476", X"0376", X"059A", X"04B0", X"019F", X"00F2", X"FFD9", X"FE28", X"016A", X"02DA", X"0767", X"0760", X"0616", X"05AC", X"00D7", X"001E", X"FDEC", X"FEDE", X"FBF4", X"FC36", X"0070", X"048D", X"0903", X"08C2", X"057D", X"0434", X"0226", X"0475", X"0199", X"022C", X"04EB", X"00F6", X"FF76", X"00C5", X"00F0", X"00DC", X"008C", X"02C4", X"06E6", X"0A75", X"0851", X"04A5", X"0101", X"FE7D", X"FF57", X"FD12", X"FDE6", X"FCB0", X"0216", X"07D4", X"090D", X"073C", X"03ED", X"0216", X"01EB", X"01E5", X"02E7", X"034E", X"043F", X"00C8", X"01C8", X"00D8", X"FF99", X"0112", X"02C5", X"04D8", X"0AC3", X"0B4A", X"0762", X"018B", X"003B", X"012E", X"FF56", X"FECE", X"FDAC", X"FDDA", X"0567", X"085D", X"0613", X"0630", X"0284", X"0229", X"028C", X"018F", X"01F1", X"0351", X"0166", X"FDF6", X"FD71", X"0009", X"FE60", X"014E", X"030F", X"038A", X"0893", X"0580", X"01B6", X"01C6", X"01F9", X"02FB", X"FF99", X"FEF6", X"FE50", X"00C3", X"048E", X"03DC", X"0447", X"03F4", X"031F", X"03DA", X"05B3", X"035D", X"01C9", X"0266", X"010B", X"FD9C", X"FD90", X"01CA", X"0045", X"0197", X"0347", X"02A0", X"0261", X"FF22", X"0196", X"00A5", X"02B7", X"0233", X"0284", X"00E5", X"0272", X"018A", X"0326", X"019E", X"0126", X"0147", X"01C9", X"053D", X"0805", X"0312", X"01C4", X"01F7", X"0175", X"FEC7", X"FF33", X"FFF1", X"0030", X"01E8", X"015F", X"FF73", X"FC56", X"FF1B", X"00C9", X"01C0", X"0360", X"0349", X"0347", X"05B0", X"0464", X"03C2", X"01AB", X"0044", X"FFCE", X"0117", X"009C", X"0393", X"0550", X"072C", X"0226", X"FEEA", X"FD90", X"FED0", X"FFC0", X"FE82", X"FFFE", X"019B", X"0018", X"FF01", X"FA0E", X"FDBD", X"FF02", X"01A0", X"0263", X"0485", X"06CB", X"05FC", X"04FF", X"0351", X"FECB", X"FDB4", X"FBD9", X"FAAB", X"FD2D", X"0355", X"0610", X"0752", X"018F", X"01D4", X"FE55", X"FD44", X"FFD4", X"00CC", X"FFB6", X"023E", X"0497", X"0101", X"FA7F", X"FAAC", X"FF32", X"FF5A", X"00D6", X"02ED", X"030A", X"01C1", X"0485", X"024A", X"FE36", X"FB76", X"F863", X"FB37", X"FE8F", X"058C", X"07D8", X"0439", X"044E", X"FDBC", X"FCD5", X"FD43", X"013F", X"FF82", X"FF9D", X"FFCC", X"02FB", X"02CB", X"FE47", X"FD5C", X"0004", X"014B", X"02FA", X"0529", X"048A", X"04F5", X"07FF", X"04C9", X"02DC", X"0470", X"FE82", X"FE47", X"FF9E", X"04B0", X"029D", X"0134", X"001A", X"FEB2", X"FD65", X"FDC3", X"FEB9", X"FF35", X"0075", X"0019", X"028B", X"0003", X"03E8", X"0478", X"057D", X"0247", X"02ED", X"0AF2", X"08AA", X"08C8", X"0851", X"0763", X"0707", X"0A36", X"07CA", X"0323", X"020D", X"00E3", X"0020", X"FFC5", X"FBF0", X"FF93", X"FEFB", X"0009", X"021F", X"0143", X"FF73", X"002F", X"004B", X"FF0C", X"02E9", X"02C9", X"03ED", X"035E", X"04F4", X"0595", X"087D", X"0999", X"07D0", X"087B", X"0639", X"0418", X"039A", X"005A", X"FFC1", X"007C", X"FFB0", X"FF71", X"00F4", X"000C", X"FFD3", X"0033", X"FFE7", X"003B", X"FFDA", X"00C3", X"FE11", X"FEE6", X"FF2A", X"FFD7", X"0050", X"01FE", X"FFD8", X"0480", X"019A", X"02DD", X"033D", X"0266", X"023B", X"006F", X"0037", X"FFF3", X"002A", X"004D", X"0138", X"012B", X"FF7A", X"0021", X"FF2C", X"00C3", X"0022"),
        (X"0082", X"FE3F", X"FFF8", X"00BA", X"0045", X"005E", X"00F6", X"FF5E", X"FEEB", X"019D", X"0048", X"0100", X"01F2", X"01FF", X"FE28", X"FE77", X"0063", X"001B", X"FF07", X"0162", X"FF1E", X"0013", X"003D", X"FFEF", X"FFE0", X"FF24", X"0027", X"FFC8", X"0117", X"0065", X"FF49", X"FF0B", X"00BB", X"008E", X"00F0", X"02FF", X"0441", X"03F4", X"04A6", X"0555", X"0551", X"056E", X"02CF", X"001C", X"FF4B", X"02CD", X"0385", X"056C", X"038D", X"03B8", X"017A", X"01BF", X"FF61", X"002E", X"0104", X"FF06", X"0035", X"00EC", X"FF7E", X"016B", X"002C", X"0102", X"0389", X"044F", X"04DC", X"0486", X"0484", X"0578", X"03BD", X"03B6", X"02F6", X"043F", X"022B", X"048A", X"060C", X"06DE", X"0867", X"07C1", X"0695", X"010C", X"FFB1", X"FE48", X"0036", X"FEB7", X"000A", X"0137", X"FEB8", X"013F", X"010D", X"FD42", X"004E", X"FDBB", X"01CB", X"FF9A", X"00A9", X"0019", X"FF45", X"0018", X"01A8", X"00D1", X"01D8", X"04C0", X"042B", X"0914", X"08BB", X"0A9E", X"083B", X"0534", X"017B", X"0041", X"00FC", X"0055", X"FF87", X"FFDA", X"FF8F", X"02B0", X"FE31", X"FC45", X"FDE8", X"FDCF", X"FA82", X"FA55", X"FC62", X"FCC9", X"FE5B", X"FA80", X"FDA4", X"FD6D", X"001D", X"0286", X"01EE", X"01ED", X"041B", X"070C", X"0746", X"0A45", X"06EF", X"018D", X"FE7B", X"FFE1", X"FE5C", X"FE94", X"FE62", X"FF4B", X"FB65", X"FCF4", X"FF9D", X"FF0A", X"FE96", X"FD40", X"FF85", X"FCC2", X"FBA6", X"FC0C", X"FCA9", X"FB15", X"FDEE", X"012D", X"0322", X"02F1", X"0270", X"0551", X"06B1", X"0736", X"04DA", X"02A7", X"0084", X"008D", X"FF02", X"FED2", X"03E6", X"0308", X"01CA", X"053D", X"FFC7", X"0162", X"0121", X"FF1D", X"FE38", X"FC4C", X"FC7B", X"FB94", X"FB30", X"F7CE", X"F74A", X"FC7D", X"FF34", X"0138", X"FFCC", X"03DC", X"0642", X"06C9", X"044E", X"00B3", X"019C", X"FF3C", X"0002", X"003E", X"01F0", X"0722", X"FFDD", X"05FE", X"04B3", X"059A", X"0386", X"038F", X"01A7", X"01D9", X"FEDE", X"FD21", X"FA4C", X"F85E", X"F9F7", X"FF03", X"014C", X"00DA", X"FF59", X"0160", X"04AC", X"042F", X"0336", X"0204", X"016F", X"FFC3", X"0018", X"05BD", X"03E6", X"04BD", X"0219", X"059E", X"056A", X"06E9", X"04BF", X"0501", X"03A6", X"0532", X"04FC", X"0047", X"F9B0", X"F836", X"FA8E", X"FEF1", X"FFCC", X"FF5C", X"012D", X"FF9C", X"FEED", X"0473", X"05FA", X"0336", X"FE82", X"FCD5", X"01A1", X"046D", X"03D4", X"0132", X"0332", X"0457", X"0255", X"0451", X"0359", X"03FB", X"0451", X"0755", X"0692", X"0423", X"FD91", X"F6E3", X"FADD", X"FD90", X"002F", X"FF67", X"FDD9", X"FED7", X"FF63", X"03E4", X"089C", X"079F", X"FFF4", X"01C6", X"0379", X"0663", X"0745", X"003F", X"01B0", X"0102", X"FD4D", X"0109", X"00B2", X"0420", X"03DC", X"03BE", X"05A9", X"0327", X"FCFC", X"F5D2", X"F9FC", X"FFAB", X"FD84", X"FDDD", X"FD69", X"FE1E", X"000D", X"014A", X"08EC", X"0840", X"0241", X"FE3E", X"0175", X"044E", X"0820", X"0267", X"FFB5", X"FD1A", X"FEC9", X"FF27", X"FF7C", X"01EE", X"03BE", X"0530", X"06C8", X"02C6", X"F4D1", X"F5C9", X"FD22", X"0030", X"FDD1", X"FBC0", X"FA4D", X"FC13", X"FEB0", X"03AC", X"03F6", X"01FA", X"FD68", X"FD36", X"FFB7", X"069A", X"09E7", X"01D5", X"FD53", X"FE8C", X"017A", X"026F", X"00FD", X"00F3", X"03F5", X"072E", X"07CB", X"FD66", X"F388", X"F66B", X"FE1E", X"FF00", X"FE0D", X"F950", X"F8D4", X"FCC4", X"0094", X"0413", X"03A7", X"FE09", X"FC53", X"FFF7", X"FFFD", X"0404", X"07F9", X"0168", X"FECC", X"006E", X"0210", X"01D8", X"0224", X"0259", X"0509", X"079A", X"03BB", X"F967", X"F607", X"F930", X"FD78", X"FDEE", X"FDB2", X"FAD2", X"FB84", X"0068", X"059F", X"0992", X"0929", X"0038", X"F88A", X"FD47", X"0198", X"040D", X"0848", X"017F", X"FFFE", X"01B9", X"035C", X"03E1", X"02BF", X"0337", X"0480", X"03B7", X"FFCB", X"F74F", X"F6D7", X"FBBD", X"FF61", X"FEE7", X"FD49", X"FDF0", X"0026", X"0562", X"0A3A", X"0C4F", X"0A45", X"FFFD", X"F84C", X"FD33", X"02A0", X"FF6C", X"0657", X"FFE9", X"FC4D", X"0078", X"0219", X"047F", X"0336", X"039B", X"0342", X"0124", X"FD1C", X"F83C", X"F85A", X"FBEB", X"FD0E", X"0068", X"FFC4", X"02A2", X"05D0", X"0AA6", X"0891", X"0B36", X"0750", X"FF63", X"FB4C", X"FE38", X"FEED", X"0191", X"0011", X"FFA1", X"FBFF", X"FE52", X"0103", X"FF8F", X"014F", X"0144", X"015D", X"0000", X"F9F2", X"F7A1", X"FB3D", X"FE46", X"FC54", X"FF43", X"01CD", X"0525", X"081B", X"076A", X"052A", X"0531", X"03B5", X"FB1C", X"F799", X"FDC5", X"00CD", X"FFA3", X"FE6A", X"FC9C", X"FF18", X"00E6", X"00FE", X"FF9B", X"FD74", X"FDAE", X"FF62", X"FE23", X"F934", X"F7F2", X"FC61", X"FD96", X"FE03", X"0057", X"04A6", X"03F7", X"053E", X"047E", X"02F0", X"0343", X"0189", X"FA98", X"F966", X"FD75", X"0072", X"0001", X"016A", X"FEDD", X"FEAB", X"012B", X"FE46", X"FDD6", X"FE92", X"FD30", X"FEDB", X"FDC5", X"FB7F", X"FD30", X"FEB8", X"FDE7", X"FFB6", X"019E", X"0353", X"041F", X"0225", X"0128", X"00B7", X"0046", X"FCE2", X"FB04", X"FA72", X"FD70", X"FFE7", X"024B", X"0207", X"FEC5", X"003A", X"FE8D", X"002A", X"FF09", X"FE9E", X"FCB6", X"FCFF", X"00AF", X"0176", X"02AA", X"016E", X"0163", X"0137", X"0203", X"0196", X"00DF", X"FEF4", X"FFAD", X"FEFB", X"FCFB", X"FDD7", X"FBF2", X"FC39", X"FDBA", X"FF28", X"FF98", X"FF72", X"FF57", X"FF11", X"FF6F", X"FD78", X"FDCD", X"FD90", X"FE3D", X"0093", X"01DB", X"059C", X"0292", X"02AE", X"0362", X"0178", X"0109", X"FFAD", X"FE0D", X"FDAD", X"FCAF", X"FC60", X"FCDA", X"FC4F", X"FAE0", X"009C", X"00CE", X"004D", X"FF40", X"FBFD", X"FD90", X"FF24", X"FDF4", X"FD58", X"FD92", X"FE22", X"FF4A", X"00E1", X"046B", X"04CA", X"045B", X"031F", X"032F", X"011C", X"00CA", X"000B", X"FE0F", X"FE6D", X"FE82", X"FD7F", X"FDFA", X"FCEE", X"FC7B", X"00CA", X"0005", X"0025", X"0043", X"FB83", X"FCD2", X"FEF2", X"FE59", X"FA95", X"FAE6", X"FC7E", X"FFF6", X"FF90", X"0205", X"0195", X"03B4", X"0223", X"0160", X"0114", X"0276", X"01E7", X"018E", X"FF17", X"FE78", X"FE7E", X"FDFF", X"FF26", X"0027", X"0338", X"FE6A", X"0115", X"019B", X"FC6D", X"FE6B", X"FFCA", X"0083", X"FE28", X"FD09", X"FEC7", X"00AD", X"0222", X"012B", X"010E", X"007C", X"02BD", X"02DC", X"01BD", X"00FD", X"FE99", X"FF70", X"FDCB", X"FD7A", X"FB79", X"FC6D", X"FE6A", X"FF79", X"00CF", X"FF9C", X"0008", X"0028", X"FFE9", X"0080", X"006F", X"0075", X"FED0", X"FF84", X"FF15", X"025A", X"01BF", X"01CD", X"01E6", X"025F", X"03E0", X"01B1", X"023C", X"00D3", X"FF15", X"FEFB", X"FB70", X"FC56", X"FBFD", X"FCD2", X"FEEB", X"FCB4", X"FE5A", X"FE32", X"FFC6", X"003B", X"FDBF", X"0111", X"022F", X"FEB1", X"FD3D", X"FD99", X"02D7", X"0277", X"005A", X"024C", X"00F8", X"FF5D", X"FF03", X"0193", X"015C", X"FE8E", X"FEB3", X"FC36", X"F9C8", X"FC4C", X"0069", X"FF6F", X"0129", X"FF11", X"FFCC", X"FF0E", X"0133", X"0106", X"FF7A", X"FF76", X"FE33", X"FDE5", X"FE68", X"0100", X"029E", X"01DB", X"004C", X"FF74", X"FF31", X"FFE2", X"FCA4", X"00B2", X"FD82", X"FDDB", X"0005", X"FFBE", X"FEDB", X"FC89", X"FE33", X"FC4C", X"FCF3", X"01B0", X"FFEE", X"00A7", X"0084", X"FF98", X"FFB6", X"002D", X"01AF", X"0234", X"00B3", X"FE2C", X"0000", X"0075", X"0081", X"FF8F", X"009D", X"06FE", X"FE4D", X"FE7B", X"0245", X"0439", X"031D", X"02B7", X"0054", X"0101", X"FE9C", X"0440", X"0009", X"0025", X"005D", X"FE57"),
        (X"FF05", X"FFE1", X"0133", X"FF4F", X"FD88", X"FF91", X"0011", X"0052", X"FF7C", X"00A8", X"FFC1", X"0040", X"FE6C", X"FECC", X"002F", X"FFBE", X"FF5C", X"FF64", X"00DF", X"0134", X"FFBA", X"FF45", X"0086", X"FF04", X"008F", X"00BF", X"0128", X"0017", X"FEE2", X"00F2", X"FECA", X"FFEA", X"FE3F", X"0030", X"0088", X"FF96", X"001F", X"0158", X"0134", X"021C", X"01FB", X"0388", X"0181", X"FE63", X"0373", X"02D1", X"0028", X"FFE0", X"0222", X"FFEC", X"0120", X"FFE8", X"0009", X"FF7F", X"FF7E", X"FEFC", X"FF08", X"FFF3", X"00FB", X"FFEA", X"FFF4", X"01E6", X"0127", X"047C", X"0548", X"0477", X"06CA", X"0546", X"0442", X"01CC", X"02EA", X"015D", X"0045", X"010C", X"00F9", X"014A", X"0049", X"03FE", X"01B4", X"0365", X"0385", X"02B3", X"FFC0", X"FE8F", X"FFDA", X"0045", X"FE9F", X"FF65", X"FEAB", X"0119", X"FEBA", X"0053", X"FF5D", X"FEE2", X"FF15", X"000D", X"FE4B", X"00A3", X"0063", X"FD8A", X"005E", X"FF6E", X"FE2F", X"FE19", X"FC3D", X"FC4B", X"FE44", X"FE38", X"FF28", X"FF81", X"01BD", X"FF76", X"FE5D", X"FE93", X"FC4E", X"FD32", X"FBB1", X"FDEB", X"FD2D", X"FE42", X"FE55", X"FE39", X"FC21", X"FC90", X"FD79", X"FDAB", X"FC07", X"FC8F", X"FE6C", X"FD84", X"FD5F", X"FCFC", X"FC73", X"FC0D", X"FCDF", X"009D", X"FE02", X"FDAC", X"FD38", X"FFCD", X"FF23", X"FF01", X"FEBC", X"FDB1", X"FF36", X"FF2E", X"FE52", X"FE3E", X"0076", X"0003", X"005B", X"FF28", X"FF84", X"FE7F", X"00AD", X"0163", X"030E", X"02A3", X"0390", X"0238", X"FF6D", X"010A", X"FFB3", X"0378", X"005F", X"FCF3", X"FF72", X"FFF7", X"0018", X"FDEF", X"FFEF", X"0038", X"0051", X"00F4", X"00AE", X"00BB", X"FE76", X"FFF1", X"FD7D", X"FE62", X"FCAC", X"FD1C", X"FF54", X"FF66", X"008E", X"0106", X"FFB3", X"0043", X"FF0A", X"FF82", X"01AF", X"01A5", X"FD76", X"FBE0", X"FDF9", X"00AF", X"FFE0", X"FC7C", X"01CF", X"FF26", X"FF7A", X"006A", X"020A", X"0060", X"FD2A", X"FEC3", X"FD06", X"FFA9", X"FD0B", X"FDE6", X"FD48", X"FDBC", X"FF3E", X"FE86", X"FDE9", X"FEF5", X"FE69", X"0096", X"01AC", X"0014", X"FCC6", X"F8D2", X"FB9A", X"FEB8", X"024D", X"00C9", X"FF51", X"FCE7", X"FF10", X"001D", X"FF9B", X"FE14", X"FE6A", X"FF3A", X"004B", X"FD93", X"FCC1", X"FE24", X"FE84", X"FFFA", X"01B1", X"01F9", X"FE70", X"FEF5", X"FF31", X"FE48", X"FD6A", X"FD6E", X"F844", X"F564", X"F9F2", X"FC85", X"FF58", X"FD24", X"FEF8", X"FC11", X"FB90", X"010F", X"FED9", X"FF51", X"FCCF", X"FFBB", X"00DB", X"FE04", X"FEA7", X"FECE", X"FF2B", X"00C9", X"0383", X"0193", X"0063", X"FF28", X"FF01", X"FDBC", X"FC6C", X"FBDD", X"F8CD", X"F3BD", X"F6D6", X"FC7D", X"FEB7", X"FDAB", X"FDE0", X"FE37", X"FC72", X"01F4", X"012E", X"FDE8", X"FBE9", X"FDC3", X"FC08", X"FD2F", X"FF2D", X"FBFF", X"FBC9", X"FE1A", X"FE99", X"00CA", X"FE93", X"FE87", X"FCDD", X"FE57", X"FB6D", X"FAC0", X"F6B0", X"F2CB", X"F4FF", X"FDA1", X"FF90", X"FDEC", X"FB9D", X"FD5F", X"FB07", X"FF37", X"0325", X"FF2F", X"FFF4", X"FD27", X"FEC2", X"FB38", X"FB84", X"F7EA", X"F585", X"F740", X"FE0D", X"FD8D", X"FDD4", X"FFE1", X"FD25", X"FF17", X"FEDC", X"FC11", X"F944", X"F40F", X"F7F2", X"FE9F", X"00B9", X"FE37", X"FCD9", X"FC83", X"FAC6", X"0009", X"0208", X"0197", X"0230", X"FE30", X"FE48", X"FD69", X"FE09", X"F967", X"F65D", X"F7B6", X"FAB3", X"F9FE", X"FD66", X"FE2F", X"FEAD", X"03A1", X"0483", X"0279", X"050E", X"FDD7", X"FD5A", X"FE04", X"FFB7", X"0174", X"FDEF", X"FB47", X"FBF4", X"FF8D", X"0324", X"0440", X"0475", X"0250", X"009D", X"FDFB", X"FC29", X"FAE6", X"F748", X"FA23", X"FA8B", X"FDDE", X"FDBD", X"FEC7", X"00DD", X"0444", X"07A6", X"0932", X"07F1", X"02FA", X"044C", X"030D", X"FFE2", X"FE19", X"FD77", X"FC99", X"FDB9", X"00AB", X"0634", X"083D", X"086E", X"05D3", X"05DA", X"02E0", X"FDB9", X"FACE", X"FA31", X"F85E", X"FBB9", X"FFE0", X"FFB6", X"00F2", X"0159", X"025E", X"0532", X"08E5", X"0978", X"06B2", X"04B3", X"0268", X"FF68", X"FDE5", X"000C", X"FE5E", X"024D", X"01AE", X"02E1", X"0621", X"080A", X"0907", X"0821", X"068D", X"01D5", X"FF6F", X"FC65", X"FCAE", X"00A1", X"0162", X"FF3D", X"0110", X"00CA", X"FF61", X"00D8", X"05C0", X"08D3", X"0B72", X"05C1", X"01F6", X"FF01", X"FDE0", X"FF5F", X"FE1B", X"FFAB", X"FEF4", X"FF77", X"02E3", X"0345", X"07E0", X"061D", X"073B", X"04EB", X"0100", X"0028", X"FF71", X"02AE", X"02AA", X"FFAD", X"00AA", X"FF99", X"0011", X"015D", X"073F", X"0E1A", X"0DBE", X"0651", X"021C", X"FFDB", X"FDBC", X"00CA", X"FC46", X"FE5D", X"FD3F", X"FE60", X"FFBD", X"0054", X"0384", X"07CE", X"0680", X"0382", X"014F", X"0097", X"0109", X"0125", X"011F", X"0109", X"FFC8", X"FF7D", X"FE67", X"0139", X"0609", X"0B5C", X"09E3", X"034A", X"04B4", X"FE1A", X"002F", X"FE14", X"FCD6", X"FE53", X"FE63", X"FC78", X"FFCB", X"0182", X"0139", X"066E", X"06EB", X"0567", X"028B", X"FF86", X"0016", X"01AC", X"FF1D", X"FF81", X"FE33", X"FD15", X"FE09", X"031F", X"0A83", X"0FD4", X"0704", X"0062", X"027C", X"FF90", X"FF13", X"FEA3", X"0131", X"FFA1", X"FE91", X"0009", X"002A", X"FE2A", X"0000", X"04B2", X"05EA", X"04CC", X"021C", X"008F", X"012A", X"009A", X"0271", X"FFCF", X"FE7E", X"FE88", X"0224", X"042A", X"05BC", X"09C5", X"0392", X"01D0", X"0063", X"FE99", X"0139", X"0173", X"0077", X"024D", X"026D", X"017C", X"007C", X"FFD1", X"FFD5", X"021E", X"051D", X"028A", X"01EA", X"0291", X"00D6", X"03E2", X"01F6", X"0378", X"01CA", X"01ED", X"02B8", X"041C", X"0795", X"09C7", X"058A", X"02D4", X"FF09", X"FFC0", X"00BF", X"02C6", X"026C", X"01CC", X"0047", X"0068", X"00A1", X"0191", X"0068", X"0227", X"027F", X"0423", X"014B", X"021E", X"039B", X"0360", X"033C", X"0467", X"030A", X"03D1", X"0380", X"075F", X"0A0C", X"081B", X"0504", X"0286", X"00A0", X"FF81", X"FEF0", X"0155", X"0180", X"008B", X"0317", X"010F", X"013F", X"024D", X"03C5", X"02E7", X"010F", X"0200", X"0053", X"FFB5", X"02DD", X"03B9", X"02B2", X"03D6", X"0279", X"0476", X"06B6", X"0900", X"0A81", X"06B6", X"02FC", X"0211", X"0185", X"0053", X"FF42", X"0029", X"FC76", X"FD7F", X"009A", X"0032", X"010C", X"02C9", X"0547", X"0215", X"0385", X"013E", X"FF91", X"0021", X"FED0", X"001A", X"01AC", X"03A7", X"02D6", X"02E0", X"04F6", X"07D4", X"0677", X"034D", X"0441", X"0177", X"FF96", X"FF9D", X"0109", X"FE7C", X"F845", X"F9E5", X"F9E7", X"FAA4", X"F88E", X"FC90", X"FD85", X"FCA6", X"FEFD", X"FEF4", X"FF6C", X"FDA3", X"FC32", X"FC9D", X"FDE5", X"FF3C", X"FD7A", X"FE74", X"00DB", X"03F7", X"04BE", X"0573", X"03E9", X"00FB", X"0181", X"00CA", X"00DE", X"019D", X"FA80", X"F9F1", X"F8C6", X"F79B", X"F406", X"F101", X"F049", X"F091", X"F021", X"EE52", X"F0C1", X"F2DE", X"F4E2", X"F478", X"F21F", X"F6DD", X"F59F", X"F635", X"F784", X"F995", X"FD03", X"FB55", X"015B", X"046E", X"FECA", X"FE83", X"005E", X"00B7", X"00BA", X"01CE", X"FFD3", X"FF3B", X"FAAC", X"FAC6", X"F60F", X"F7C1", X"F752", X"FB02", X"F56B", X"F283", X"F466", X"F32D", X"F33F", X"F557", X"F699", X"F57E", X"F587", X"FA28", X"FE7D", X"FE74", X"01BB", X"FFAD", X"00B2", X"FF96", X"009A", X"01D5", X"FFDC", X"0012", X"0084", X"FD4C", X"FCC5", X"FB79", X"FBD3", X"FBA9", X"FCAE", X"FCCC", X"FC1C", X"FAD9", X"FB24", X"FCE1", X"FD17", X"FDC2", X"FE2D", X"FC98", X"FC6E", X"FA88", X"FB7E", X"FFEB", X"009B", X"00AC", X"0070"),
        (X"FFD1", X"00B0", X"00E9", X"FF20", X"00C4", X"FFA8", X"0051", X"FE8A", X"0041", X"0014", X"006F", X"0007", X"FE99", X"FEF0", X"002E", X"007F", X"FED3", X"FF97", X"FF92", X"FE9F", X"00C2", X"001F", X"FEBB", X"00DE", X"0054", X"FECB", X"FFF0", X"010E", X"00BB", X"FFDA", X"FE64", X"FEE7", X"009E", X"0043", X"FF8B", X"FE26", X"FBA4", X"FC31", X"FD67", X"FC01", X"FBFF", X"FB84", X"0002", X"00A0", X"02F2", X"FF99", X"FB95", X"FC58", X"FC2A", X"FDED", X"FCD4", X"FF93", X"FFCD", X"FFD8", X"FFC5", X"FFCB", X"004C", X"FF61", X"FEDB", X"011E", X"FE07", X"FE38", X"FEEC", X"FC7E", X"FD07", X"FE2C", X"FC6C", X"FD82", X"FE9D", X"FEF4", X"FF5F", X"0331", X"028B", X"00B0", X"003E", X"FDE6", X"FD4D", X"F9E4", X"FB25", X"FC29", X"0117", X"0227", X"007A", X"FF7A", X"008D", X"0022", X"000E", X"FF4D", X"01D4", X"FE6F", X"FD41", X"FE26", X"FEA0", X"FEA8", X"FF96", X"FF23", X"017A", X"0317", X"049B", X"0469", X"03B0", X"045B", X"043F", X"00CC", X"00EB", X"FDF4", X"FDCE", X"FBB1", X"FEED", X"0009", X"FE6D", X"FF43", X"FFEC", X"FF9D", X"FFDE", X"00F6", X"FCEA", X"FCF5", X"0288", X"FFBB", X"FF9A", X"01C1", X"032B", X"0444", X"04A1", X"FFFF", X"01AD", X"03BC", X"02F9", X"026C", X"02FD", X"FEDD", X"FEF7", X"FDFA", X"FD9D", X"FDBB", X"01EB", X"01EF", X"01DD", X"FE6B", X"0049", X"003C", X"0141", X"01DD", X"FD85", X"FE36", X"FD36", X"FFFA", X"00C8", X"0314", X"0293", X"05D4", X"0400", X"04EB", X"01F3", X"018E", X"0220", X"012F", X"FF04", X"FE92", X"00A8", X"00C9", X"FDEC", X"FED0", X"0058", X"0376", X"00D4", X"FD73", X"01A7", X"FE80", X"FF46", X"01E5", X"FFC3", X"FE8D", X"FBF8", X"FE9A", X"FF94", X"021D", X"0404", X"048D", X"04A2", X"06FB", X"05EF", X"06B0", X"0649", X"048C", X"0444", X"0418", X"01B2", X"FDEA", X"FCB8", X"FE09", X"0217", X"0507", X"05A6", X"FFDD", X"004E", X"FF1F", X"01F1", X"01B9", X"FEAF", X"FDE2", X"011D", X"FE28", X"0115", X"00E0", X"0218", X"02E4", X"03E2", X"038D", X"03EE", X"04F9", X"041C", X"03A6", X"02E8", X"038F", X"01D1", X"FF39", X"FF95", X"FE65", X"00F9", X"0677", X"0332", X"0031", X"FE71", X"FED0", X"FE49", X"FE3D", X"FAB4", X"00DF", X"017C", X"0077", X"02B1", X"0056", X"0287", X"0344", X"022A", X"0433", X"0401", X"03CF", X"011E", X"0118", X"01B3", X"0187", X"00E0", X"0282", X"0176", X"0087", X"0668", X"0A67", X"07E4", X"04C5", X"0033", X"FE5C", X"006C", X"00E9", X"FDEA", X"0323", X"04D8", X"0441", X"0049", X"0236", X"0229", X"038F", X"0303", X"0283", X"03D3", X"05C3", X"FF93", X"00A0", X"0043", X"FF61", X"013F", X"0190", X"015C", X"016F", X"0872", X"0EFF", X"0B14", X"0234", X"010E", X"FFC1", X"FE64", X"0110", X"FF5C", X"0323", X"05F7", X"022D", X"00AD", X"FFC4", X"00EE", X"FFCD", X"FE75", X"FE81", X"0608", X"058F", X"00E0", X"FE33", X"FF9D", X"FF20", X"FE44", X"00A1", X"FFC8", X"0088", X"069F", X"0DED", X"0AD2", X"02AD", X"FFF0", X"FCFE", X"FDB1", X"FE84", X"00EF", X"0228", X"03B0", X"00D2", X"FE6D", X"FDFB", X"FE5B", X"FC42", X"FB03", X"FCB1", X"063A", X"04C7", X"FF08", X"FE5A", X"FF4B", X"FEB3", X"FE59", X"FC76", X"FB8F", X"FC90", X"FE19", X"0B1B", X"0ACE", X"0277", X"FFAA", X"FF01", X"FECE", X"FE45", X"05FA", X"0283", X"FE0C", X"FE03", X"FBCF", X"FA6D", X"FA30", X"F9FE", X"F8E2", X"FF2A", X"06F3", X"03DB", X"FE41", X"FE15", X"FF1A", X"FF90", X"FEEC", X"FCB9", X"F837", X"F700", X"F679", X"01F3", X"074F", X"04FE", X"0060", X"FEC2", X"FE4E", X"FF9B", X"05EE", X"FD5D", X"FA14", X"FDBB", X"FC03", X"FB6A", X"FB2D", X"F974", X"FA7C", X"05A6", X"07C6", X"029B", X"FF51", X"FF04", X"FED7", X"006B", X"00E8", X"FE80", X"FA51", X"F5D0", X"F9B8", X"025D", X"07A9", X"0193", X"0188", X"0109", X"FEF9", X"009C", X"037C", X"FC8D", X"FBE3", X"FB7F", X"FB3B", X"F92A", X"F95E", X"F812", X"FCF2", X"070D", X"077F", X"0497", X"FFE5", X"00EA", X"0146", X"FFAB", X"FF14", X"FEAE", X"FC94", X"FA39", X"FCBD", X"017E", X"0793", X"02B1", X"008A", X"FF9A", X"FC2C", X"005F", X"0419", X"FE27", X"FC23", X"FDA4", X"F94F", X"F90A", X"FA06", X"FA57", X"FEE0", X"05D9", X"03F2", X"02EB", X"00B3", X"FFCC", X"FFFC", X"0087", X"01A5", X"FEFE", X"FCFB", X"FD4A", X"0060", X"028C", X"0798", X"02DA", X"FF09", X"FFC0", X"0113", X"05FF", X"0767", X"0274", X"FE73", X"FBFB", X"FC3F", X"FA7D", X"FD84", X"FC10", X"01B3", X"04F7", X"03C8", X"0103", X"0006", X"0065", X"FF46", X"FD9F", X"FE52", X"FDA2", X"011E", X"00CD", X"01AE", X"0361", X"06C8", X"0356", X"FF87", X"FEF0", X"FEEE", X"068E", X"04ED", X"037D", X"03C8", X"FFF1", X"FD87", X"FE57", X"FC7E", X"FCA9", X"013F", X"03BB", X"02D7", X"0231", X"FF6C", X"FE43", X"FE3A", X"0131", X"FDCB", X"FEE2", X"0106", X"02C5", X"032A", X"0526", X"07F8", X"024F", X"02F2", X"0144", X"FEA2", X"0344", X"0479", X"0634", X"0580", X"00CB", X"FF0F", X"FDE8", X"FF15", X"FEDA", X"FF67", X"0250", X"0377", X"02A9", X"FF9C", X"FF70", X"FECA", X"FF86", X"0009", X"FF90", X"016E", X"026B", X"04B6", X"0540", X"04AF", X"04EC", X"FF07", X"FC6C", X"FED2", X"024D", X"01A4", X"0257", X"03F6", X"038C", X"FF76", X"FDCB", X"FEC3", X"FC81", X"FE72", X"0139", X"00E3", X"FF56", X"FF15", X"FF7D", X"0009", X"0079", X"FF72", X"FD90", X"03F7", X"059D", X"061E", X"076D", X"042B", X"01FC", X"0201", X"FD32", X"FEC8", X"023A", X"00D6", X"024D", X"03CF", X"0369", X"019C", X"FE0D", X"FD04", X"FDC5", X"FC06", X"FE8A", X"FC56", X"FD8F", X"FE5B", X"00D9", X"FDD3", X"009E", X"FFF1", X"00D3", X"074A", X"0713", X"08A1", X"07BF", X"012B", X"0118", X"FFCE", X"007E", X"01D2", X"014C", X"02BF", X"FFDB", X"0457", X"0326", X"0141", X"0018", X"FE20", X"FB35", X"FBB4", X"FD1F", X"FC29", X"FCFA", X"FF6A", X"0034", X"FFB5", X"00D6", X"008A", X"0275", X"0420", X"05DA", X"0624", X"05F8", X"FD82", X"FF92", X"FF50", X"00A3", X"00CD", X"0436", X"0435", X"FFD0", X"0008", X"028C", X"0162", X"0141", X"FE10", X"FCB9", X"FDD5", X"FD99", X"FF69", X"FCC2", X"0102", X"00E6", X"0087", X"FEE7", X"0164", X"FF14", X"0194", X"056F", X"0465", X"03B8", X"FD96", X"FFE4", X"FFA6", X"FF55", X"0122", X"04A1", X"0538", X"FFD3", X"FE13", X"FE21", X"FF0B", X"FEBD", X"01D4", X"FDAA", X"FFC7", X"FF3C", X"01B1", X"003F", X"FF47", X"FFDE", X"FED3", X"FEB2", X"FED9", X"FEA3", X"029F", X"04C9", X"0629", X"02CB", X"FE03", X"01D6", X"000C", X"FFC9", X"FE63", X"FEAC", X"035D", X"04DF", X"04B8", X"0682", X"038C", X"055B", X"0527", X"042C", X"0677", X"07AF", X"04ED", X"04B5", X"0250", X"0443", X"020A", X"01FA", X"04E9", X"02C5", X"0047", X"0470", X"0450", X"FED6", X"00D5", X"FF65", X"0005", X"001E", X"00A8", X"0037", X"0430", X"07C8", X"063C", X"08C8", X"0B2C", X"0B10", X"092E", X"08DC", X"09A4", X"07A3", X"06FB", X"0460", X"0479", X"04D3", X"05BB", X"05B7", X"09BE", X"07C5", X"05FC", X"04B5", X"048C", X"0162", X"012A", X"00F7", X"FFC6", X"0070", X"FEDA", X"017E", X"0376", X"0518", X"0890", X"08FA", X"08BC", X"0C07", X"0BD4", X"0C88", X"0A66", X"0B31", X"0DAE", X"0A25", X"08ED", X"081B", X"0A22", X"08A1", X"0BBB", X"08A9", X"0530", X"0297", X"01CD", X"001A", X"009F", X"00DA", X"FEA3", X"FFFA", X"01F7", X"0125", X"FFC1", X"FED3", X"031D", X"0349", X"03DC", X"0637", X"04F4", X"05D6", X"071D", X"061D", X"081F", X"06EF", X"0553", X"02C7", X"0714", X"0450", X"FF1A", X"FF51", X"005E", X"FF75", X"FF35", X"FFBE", X"004C", X"0078"),
        (X"0127", X"0002", X"0015", X"FFBD", X"0069", X"FF45", X"FE21", X"01A2", X"00D0", X"007E", X"FF7A", X"FF91", X"FE7C", X"FF81", X"FF0D", X"FFDB", X"00BE", X"00D5", X"0148", X"FF93", X"0274", X"FFCB", X"0002", X"FF59", X"00DF", X"FFD7", X"FE13", X"FEEF", X"FFEB", X"FF89", X"00B8", X"003A", X"FF78", X"00AA", X"FE8E", X"FFA5", X"FFA2", X"0147", X"FE96", X"004E", X"FF9B", X"FE35", X"02C1", X"021F", X"FCC7", X"FC06", X"FE53", X"FD45", X"FAFC", X"FCB0", X"FCB5", X"FD4F", X"FFA8", X"0208", X"00EB", X"00B1", X"FFB6", X"FF3C", X"00CD", X"FEE2", X"0009", X"FEE2", X"FF8B", X"FD36", X"FB41", X"F772", X"F774", X"F9E0", X"FBD7", X"FBB0", X"FD58", X"FE98", X"FF75", X"FE87", X"FFD3", X"FF7B", X"FC9C", X"FCA4", X"FDB6", X"FAE5", X"FC58", X"FC88", X"00FA", X"FEEE", X"FE98", X"00AA", X"0273", X"FF77", X"0101", X"FD5C", X"F8D5", X"F938", X"F786", X"F8B6", X"FB08", X"F691", X"F8F6", X"FC8E", X"FC5D", X"FED0", X"FC34", X"FDD9", X"FD47", X"FF67", X"FD89", X"FE63", X"00CF", X"0056", X"FEFB", X"FDF2", X"00DE", X"0140", X"FFE4", X"004C", X"01B1", X"FD74", X"0056", X"FC56", X"FB5F", X"FC40", X"FD94", X"0024", X"FF9A", X"FFE8", X"0296", X"041A", X"05D0", X"0838", X"048A", X"0588", X"044C", X"04DE", X"0636", X"08D3", X"0716", X"05EC", X"01E5", X"FF5F", X"FFE7", X"FFD6", X"001D", X"FFC1", X"0202", X"FDE2", X"FC6A", X"FD11", X"FDFB", X"FDB0", X"FD41", X"FEAF", X"0017", X"FF35", X"033A", X"03B2", X"05A5", X"0403", X"0450", X"04D3", X"043E", X"04ED", X"05EE", X"0934", X"0990", X"091E", X"068C", X"027D", X"02B5", X"FF1C", X"0040", X"FF39", X"FDC5", X"F9AF", X"F9B6", X"FD8E", X"0101", X"FE8C", X"FE60", X"FCF7", X"FD92", X"FEF5", X"FF68", X"FCBC", X"FB02", X"FC07", X"FD98", X"FF1C", X"FF8C", X"0495", X"067F", X"0578", X"094F", X"0CA0", X"0A96", X"06DB", X"036B", X"0250", X"005D", X"FC9F", X"FB37", X"F96A", X"FA40", X"FEC9", X"FE73", X"01A5", X"FF75", X"FD17", X"FFD2", X"FCF2", X"FB5D", X"FAAB", X"F8C9", X"FB88", X"FAE3", X"005B", X"017D", X"03CF", X"0353", X"0300", X"05FA", X"0BA8", X"0DDF", X"061F", X"0484", X"0286", X"01A9", X"FCDC", X"FD72", X"FC66", X"FB54", X"FFC3", X"FF7A", X"FE65", X"FC7B", X"FE05", X"FBA6", X"FCDE", X"FE78", X"FE62", X"FA87", X"FBB7", X"FF5E", X"0377", X"0458", X"02E8", X"0449", X"033D", X"03A6", X"0764", X"0E54", X"0B3F", X"048F", X"0223", X"FFDA", X"FB7D", X"FD83", X"FC51", X"FC66", X"FE17", X"FE38", X"FD68", X"FADA", X"FB05", X"FAC4", X"FD8F", X"FE60", X"FDE7", X"FC5E", X"FCBF", X"0064", X"030C", X"0303", X"033F", X"01AB", X"043B", X"022A", X"0590", X"0B23", X"073E", X"0420", X"FE63", X"0020", X"FEFB", X"FB1C", X"F982", X"002B", X"FD58", X"FA27", X"FCD8", X"FE87", X"FDE3", X"005A", X"0421", X"0344", X"037F", X"027C", X"02CD", X"0027", X"FDB2", X"FF93", X"FF4F", X"FFD2", X"0279", X"02B5", X"041B", X"04CC", X"04FB", X"0306", X"FF46", X"FFD8", X"FC61", X"FB96", X"FB50", X"FCAB", X"FEA8", X"FEF8", X"0110", X"01C1", X"049A", X"0791", X"066D", X"063A", X"049F", X"0354", X"0124", X"FD23", X"FC23", X"FA64", X"FB57", X"FE43", X"019C", X"022A", X"049E", X"0672", X"044F", X"05E4", X"0292", X"FF44", X"FD4A", X"FD0F", X"FE46", X"FF43", X"022A", X"0372", X"04B2", X"060E", X"0888", X"067C", X"060B", X"03DD", X"0201", X"004D", X"FEFE", X"FDF5", X"FA4D", X"FC21", X"FD50", X"FE95", X"02DF", X"0450", X"03F8", X"005B", X"FECF", X"0073", X"FE93", X"0105", X"00EF", X"FE7F", X"FFC4", X"0147", X"0437", X"045F", X"079A", X"06BA", X"0727", X"0356", X"0261", X"008A", X"FDE7", X"FDFD", X"005D", X"FD9A", X"FBD4", X"FC34", X"FE94", X"0102", X"0208", X"04DF", X"00DA", X"FCBB", X"FAB9", X"F9C7", X"FD47", X"02D1", X"0009", X"FF62", X"FE28", X"0166", X"05E2", X"04CD", X"05B4", X"0698", X"04E5", X"007A", X"FD0F", X"FD5A", X"FEA0", X"0136", X"FF29", X"FD99", X"FC98", X"FAF0", X"FD6D", X"FD83", X"012B", X"0126", X"FFFF", X"FE26", X"F8F1", X"F7D9", X"FE8E", X"01A9", X"FECC", X"0358", X"FE43", X"01C0", X"0206", X"02A9", X"03EF", X"0594", X"03D8", X"FBEE", X"FCEB", X"FCF7", X"FFD8", X"03A9", X"FFFC", X"FCCF", X"FC10", X"FBB7", X"FC77", X"FD25", X"FE79", X"FF4D", X"FF44", X"FA7E", X"F9BA", X"FAC6", X"FC4E", X"FFBF", X"FEDF", X"FD54", X"FD92", X"FD6A", X"01C1", X"0244", X"02F4", X"0286", X"0065", X"FCE8", X"FB41", X"FF29", X"0385", X"03E0", X"FEB6", X"FC7A", X"FD24", X"FC61", X"FD85", X"0050", X"FDC0", X"FDC0", X"FE7C", X"FB13", X"F671", X"F6B3", X"FD0A", X"0029", X"001C", X"FC7A", X"FB01", X"FB4B", X"012A", X"00D9", X"0354", X"03DC", X"0177", X"FF5B", X"FF70", X"FFDF", X"0128", X"FFBA", X"FDE4", X"FE46", X"FCD0", X"FCC0", X"FF28", X"FFCF", X"FE65", X"FDFE", X"FEC6", X"FC1E", X"F70D", X"F955", X"FCE8", X"FD9E", X"FFE7", X"FC4C", X"F95A", X"F9EC", X"FE43", X"0089", X"02AA", X"048B", X"0356", X"FF69", X"FEC4", X"FFEA", X"FE6F", X"FEE5", X"FE26", X"FD15", X"FD5D", X"FDE2", X"FE34", X"00F6", X"FE23", X"FEC9", X"FD01", X"FC5C", X"F813", X"FA59", X"FE4D", X"FF70", X"FD7C", X"0031", X"FA11", X"FA3B", X"FCC5", X"022E", X"0408", X"03C4", X"0483", X"01E0", X"FF62", X"FF26", X"FFE6", X"FF3C", X"FEB5", X"FF8C", X"FF5E", X"00F7", X"015F", X"0081", X"FFED", X"FF13", X"FDD9", X"FE31", X"FC8C", X"FC25", X"FFD8", X"003B", X"01AD", X"FEA0", X"F923", X"FB28", X"FC80", X"0269", X"03BC", X"0446", X"04D2", X"04F2", X"0367", X"005B", X"FF87", X"FF43", X"01B3", X"0116", X"018F", X"0194", X"00B4", X"01BF", X"00FC", X"019D", X"0004", X"FD36", X"FB63", X"FD97", X"0039", X"00A2", X"FF5E", X"F81E", X"F97B", X"FE1A", X"01DC", X"049B", X"034F", X"05B3", X"04CC", X"04B5", X"0240", X"02D5", X"033A", X"0434", X"054D", X"02F1", X"052E", X"03F0", X"02AC", X"039B", X"0329", X"0308", X"00CF", X"FBBD", X"FD07", X"0079", X"FF1F", X"015D", X"0081", X"F8C7", X"FB58", X"FCD2", X"01E7", X"0107", X"0120", X"0230", X"02C6", X"0283", X"0286", X"03CB", X"0356", X"065E", X"049D", X"04DD", X"0630", X"05A3", X"0760", X"073F", X"054E", X"0136", X"FE47", X"FCE2", X"FD78", X"04A8", X"003A", X"0034", X"01F7", X"FE3D", X"FBCD", X"FC73", X"FD20", X"FC34", X"FC5B", X"0033", X"03B7", X"0240", X"0251", X"029D", X"04D9", X"0392", X"0667", X"07EA", X"084B", X"060E", X"05FF", X"0501", X"02EB", X"FEA9", X"FC5F", X"FA66", X"FDFA", X"029E", X"001F", X"FE9B", X"FFF6", X"FEC3", X"FD96", X"F7EF", X"F918", X"F97B", X"F79B", X"FC20", X"FF8F", X"FE62", X"FE77", X"01E4", X"0150", X"023E", X"0499", X"03A7", X"0129", X"050C", X"030D", X"0017", X"FC38", X"FC4B", X"FF05", X"FBE3", X"FCAC", X"FCEC", X"FF9F", X"0072", X"0012", X"FF59", X"00DD", X"F92C", X"F63A", X"F825", X"F7D2", X"F839", X"FC54", X"FB70", X"FDCB", X"F948", X"FB23", X"FB51", X"FFB0", X"FE4E", X"FECD", X"FC9D", X"FD20", X"FA55", X"FD9F", X"0002", X"01DB", X"01BB", X"FE13", X"0030", X"009A", X"000D", X"0159", X"FFF5", X"FF2C", X"FAEC", X"FA08", X"F73D", X"F721", X"F692", X"F6E8", X"F6A1", X"F936", X"F888", X"F6B7", X"F6CA", X"F800", X"F61E", X"F5CF", X"F84F", X"F7F7", X"FAE2", X"FD78", X"FD1C", X"FDB9", X"FC82", X"FFEC", X"FE84", X"0015", X"0121", X"FF8F", X"00DB", X"00A0", X"FF32", X"01DD", X"FD87", X"FCE2", X"FB29", X"FC98", X"FA4C", X"F982", X"FBED", X"F9CE", X"F757", X"FA83", X"FA0D", X"FA08", X"F9E3", X"FB97", X"FC6C", X"FBAE", X"FCE9", X"FE04", X"FF03", X"FF83", X"0003", X"0051"),
        (X"FF11", X"00C2", X"FF75", X"0121", X"FFD7", X"FF54", X"0121", X"FF35", X"FFFA", X"FF7A", X"003C", X"0096", X"0179", X"01A1", X"0031", X"FFCB", X"FFDC", X"FE75", X"00DA", X"002F", X"0039", X"FF7A", X"FF13", X"FF7B", X"FEC6", X"0045", X"00B2", X"0044", X"FFE1", X"0159", X"FF63", X"0073", X"FF6B", X"012F", X"0351", X"03F5", X"041F", X"066D", X"074B", X"07A2", X"0907", X"0980", X"0451", X"0717", X"0424", X"05FB", X"05C5", X"061E", X"0519", X"0216", X"02FF", X"0219", X"008C", X"00BD", X"FF22", X"FFAD", X"FFA5", X"FF6C", X"00E0", X"00CD", X"0327", X"026B", X"06A2", X"077E", X"0A4F", X"0AA9", X"0CA2", X"0B2C", X"0C5A", X"09BC", X"0695", X"0773", X"056D", X"061F", X"083C", X"0812", X"080F", X"0591", X"0782", X"0511", X"FE72", X"FDAD", X"013F", X"FFA4", X"0162", X"FF69", X"FF4C", X"0273", X"0492", X"04E5", X"0553", X"059B", X"0675", X"0851", X"06E4", X"078B", X"0A6B", X"06D6", X"05F2", X"0473", X"0368", X"0396", X"0480", X"06BD", X"084F", X"0602", X"04F4", X"0412", X"00E1", X"FF05", X"0211", X"FF40", X"0080", X"0115", X"FEA6", X"03EF", X"01C4", X"0332", X"0277", X"001F", X"02C4", X"0279", X"0177", X"01F1", X"00FE", X"00E9", X"FF19", X"0281", X"0258", X"03D5", X"036D", X"013A", X"FFCF", X"00B3", X"0238", X"0347", X"FFBD", X"FF93", X"FF23", X"FEB8", X"0072", X"0020", X"FE5F", X"0103", X"FD4A", X"FF1A", X"008A", X"0059", X"023F", X"00EB", X"03AE", X"0254", X"00B0", X"00D6", X"FFA5", X"FEE8", X"FF06", X"FF26", X"FF43", X"FF14", X"FFA0", X"0009", X"FFC4", X"01D6", X"00BA", X"FF7E", X"034F", X"0096", X"FEB2", X"FF1E", X"0282", X"FE87", X"FDC9", X"FC6C", X"FD7B", X"01A2", X"00EC", X"FEE0", X"0029", X"0029", X"01E8", X"0137", X"02EC", X"0369", X"0342", X"036B", X"0273", X"FF8D", X"FDB7", X"FFB7", X"FDA3", X"FE95", X"0131", X"0283", X"01BE", X"FD6B", X"0123", X"FEB4", X"FD91", X"FEB3", X"F943", X"FB25", X"FB93", X"FE7B", X"FD81", X"FF69", X"00D1", X"0111", X"0254", X"015B", X"0506", X"06E0", X"0622", X"04E9", X"005C", X"FD99", X"FF3D", X"FD70", X"FBC3", X"FB76", X"FFB3", X"01E3", X"FFAF", X"FFA7", X"0345", X"0195", X"00BE", X"FCCF", X"F81A", X"FB05", X"FC23", X"FADD", X"FEAF", X"FD30", X"FEC5", X"FFD8", X"FFCE", X"000F", X"058B", X"083C", X"0658", X"005B", X"FC55", X"FB96", X"FCAA", X"FC13", X"F91E", X"FBB4", X"02B1", X"0243", X"007B", X"FDE0", X"0051", X"0382", X"01D8", X"0040", X"FC95", X"FB45", X"FD1A", X"FD75", X"FF7B", X"FFE1", X"0099", X"0060", X"0271", X"0405", X"0A5C", X"06DC", X"FF72", X"F989", X"FA25", X"F9C8", X"FA5C", X"F9BF", X"F8C0", X"FCA3", X"0411", X"05BE", X"02AF", X"0392", X"0025", X"0291", X"0405", X"021F", X"FE41", X"FC8A", X"005F", X"016B", X"0015", X"02A8", X"0341", X"0477", X"0515", X"0A0C", X"0B1A", X"00E3", X"F7A6", X"F7FE", X"FB76", X"F9B2", X"FA33", X"F929", X"F9F7", X"00CB", X"0527", X"0743", X"059E", X"FEC5", X"FFA5", X"0241", X"07B2", X"035C", X"0182", X"FFA0", X"0303", X"01F3", X"01FE", X"02B0", X"050F", X"048E", X"0355", X"04C9", X"011A", X"FA9D", X"F6D3", X"FBED", X"FEE0", X"FC20", X"FB07", X"FC86", X"FE4D", X"03FE", X"0301", X"01CA", X"FF38", X"FE33", X"FEEA", X"035E", X"05D1", X"039E", X"044E", X"0309", X"076D", X"0733", X"056C", X"03B9", X"04F8", X"0242", X"FF4A", X"FFC4", X"FCF7", X"FA7C", X"F93A", X"FDBC", X"0010", X"FBE1", X"FC0B", X"FDFB", X"009B", X"034C", X"FF60", X"FCA6", X"FECD", X"FF5F", X"01A5", X"0113", X"04C4", X"055A", X"0642", X"065C", X"068A", X"05C8", X"05E3", X"030E", X"010D", X"FE6F", X"FCFA", X"FC7C", X"FCB0", X"F9ED", X"FBD3", X"FEB6", X"FE61", X"FEB0", X"FC98", X"FF00", X"03A5", X"060E", X"01CB", X"FCBF", X"F8EF", X"FD9E", X"0175", X"008F", X"0231", X"020D", X"03B3", X"05A5", X"04E9", X"0490", X"02AC", X"01CC", X"03BD", X"FC12", X"FC12", X"FBB6", X"FC1D", X"FC09", X"FB9E", X"FCD1", X"FED7", X"FF43", X"FF34", X"03AF", X"04B1", X"0611", X"02DA", X"FA1C", X"FA0D", X"FD60", X"0116", X"00AB", X"FE28", X"FC72", X"FFD1", X"02FA", X"0064", X"004C", X"011E", X"01A4", X"023B", X"FF49", X"FF41", X"FAD0", X"FBCE", X"F9FA", X"FAD9", X"FE01", X"FF9A", X"000D", X"00F9", X"0145", X"010D", X"0312", X"0335", X"FDE8", X"F994", X"FDF2", X"FF4C", X"0275", X"FFD1", X"FD5A", X"FE63", X"FEEF", X"FBF2", X"FCE1", X"FD3E", X"014D", X"01CB", X"0300", X"FD26", X"FAAC", X"FA7D", X"F93A", X"FB1C", X"FD0D", X"0153", X"00D8", X"0015", X"FD39", X"0027", X"0063", X"FFB5", X"FDD5", X"F72E", X"FE30", X"FE85", X"0213", X"FE01", X"FEA1", X"FB9C", X"FBE1", X"FC3A", X"FAC2", X"FBE9", X"FCE7", X"FFCD", X"FDF3", X"F83E", X"F6B6", X"F9D2", X"FA48", X"FC16", X"FF22", X"0076", X"011D", X"013C", X"01A5", X"0158", X"00B7", X"FCED", X"FE82", X"FC01", X"00EF", X"03C0", X"01B5", X"021F", X"FF64", X"FE26", X"FA59", X"FC56", X"FCDE", X"FC86", X"FB22", X"FCCC", X"F9B0", X"F6D1", X"F7DC", X"FC06", X"FEE6", X"0068", X"0244", X"02B6", X"01F7", X"01AD", X"02AB", X"025F", X"FEB2", X"FC6C", X"FD5C", X"FEA2", X"FE59", X"FF42", X"04E8", X"0376", X"0017", X"FF63", X"FC5F", X"FD6D", X"FBCF", X"FE10", X"FAE1", X"FC63", X"FE26", X"00DE", X"01A8", X"0438", X"00D5", X"0182", X"01DC", X"017E", X"0319", X"0355", X"0277", X"0060", X"FF23", X"0006", X"FFF2", X"FD05", X"FF3E", X"00BB", X"037E", X"0208", X"FF9E", X"FC64", X"00B3", X"FE06", X"FE7E", X"FD2F", X"FC7A", X"FF7E", X"0059", X"04E6", X"07AD", X"05ED", X"02A8", X"00F6", X"0162", X"0058", X"0095", X"00AE", X"01CA", X"013D", X"007A", X"0163", X"02F3", X"020D", X"FF8B", X"00EF", X"FFBD", X"FEA9", X"0118", X"FF1B", X"FEFF", X"FD70", X"FDCA", X"FD66", X"FE61", X"01A9", X"0270", X"0594", X"0478", X"0279", X"0244", X"001A", X"FFD9", X"FCA6", X"FE88", X"0170", X"00D4", X"0163", X"0200", X"00FD", X"032A", X"01FE", X"0003", X"00B7", X"00D7", X"FF0A", X"0071", X"FE15", X"FE1D", X"FB38", X"FCB5", X"FD11", X"FFB2", X"0251", X"037B", X"0394", X"036E", X"005C", X"0146", X"026B", X"0021", X"FE24", X"FDB9", X"FF4F", X"FDCD", X"0194", X"0262", X"FFD3", X"02A4", X"0340", X"012D", X"0095", X"001F", X"0175", X"0361", X"00CB", X"00E5", X"FC2F", X"FA51", X"FE4C", X"0113", X"05B6", X"0402", X"0266", X"0127", X"033A", X"0170", X"FF14", X"FFE0", X"FC27", X"FA65", X"FD03", X"FE0C", X"02ED", X"03A8", X"0199", X"00A0", X"0279", X"0010", X"0049", X"000F", X"0265", X"02EF", X"01C2", X"0419", X"024E", X"0257", X"0321", X"0583", X"0394", X"01C1", X"0152", X"FEA6", X"FFED", X"FFE7", X"FF20", X"FFCD", X"FDCF", X"FE68", X"0025", X"00CF", X"03F8", X"04A5", X"02C1", X"FDB8", X"FD83", X"012E", X"FFF9", X"009B", X"01D4", X"033F", X"0114", X"0695", X"03A7", X"051E", X"08F0", X"086C", X"04FF", X"066D", X"07DF", X"0527", X"05D0", X"04A6", X"0603", X"0930", X"08EF", X"09F8", X"094E", X"0BE3", X"0819", X"075B", X"053B", X"0102", X"FD64", X"01D9", X"FF3C", X"0040", X"002B", X"019B", X"038C", X"0445", X"04A3", X"086E", X"0ACF", X"09A3", X"0949", X"0AE9", X"0E02", X"0F5C", X"1344", X"10CC", X"1078", X"0E36", X"0D7D", X"0E21", X"0DFC", X"0C8F", X"068E", X"03FE", X"017E", X"00DD", X"00C2", X"FE60", X"001F", X"0028", X"002E", X"004E", X"00C3", X"0084", X"0460", X"03DB", X"048F", X"07B0", X"06BC", X"0780", X"0779", X"0608", X"087C", X"0677", X"05F0", X"05C3", X"03FD", X"036A", X"03FB", X"03A8", X"FE0B", X"FC3C", X"00EB", X"FFB3", X"FECE", X"FF62"),
        (X"FF40", X"0095", X"009A", X"0181", X"FEEA", X"0014", X"FF97", X"FFF5", X"FFCB", X"FF11", X"FFA1", X"FFB6", X"FE75", X"FCC6", X"FFCD", X"00D8", X"0050", X"01D3", X"00B9", X"0024", X"FF13", X"00B1", X"011A", X"002E", X"008E", X"000B", X"005B", X"FFDD", X"FF6F", X"FFB1", X"FF19", X"FFBA", X"00B6", X"FFC4", X"FCAA", X"FAE6", X"FC3B", X"FB9F", X"FC39", X"F971", X"FA0E", X"F9EE", X"FDDC", X"FB29", X"FBA0", X"F964", X"FA9B", X"FAB9", X"FA9F", X"FC2C", X"FBDA", X"FD3D", X"0083", X"FF2F", X"FFCB", X"0087", X"0095", X"FFE9", X"00E6", X"FE6E", X"FCBF", X"FECD", X"FC1C", X"FAC1", X"F93E", X"F762", X"F5DA", X"F6DE", X"F5CA", X"F9BC", X"F86F", X"F573", X"F880", X"FB93", X"F802", X"FAD1", X"F789", X"F75E", X"F99A", X"F710", X"FB63", X"FD8D", X"FF70", X"FF9C", X"FF31", X"00D9", X"FFA4", X"FDD7", X"FE7E", X"FDBB", X"FBFC", X"F78C", X"F770", X"F794", X"F93D", X"FA48", X"F803", X"F550", X"F773", X"FA76", X"F95E", X"FAC2", X"FADF", X"FA96", X"F810", X"F93A", X"F940", X"F84A", X"F865", X"FB4D", X"FE65", X"007C", X"FFFF", X"FE9F", X"FD90", X"FFFA", X"FD6B", X"FD3E", X"FC6A", X"FCCC", X"F8EE", X"F8CA", X"F99F", X"F898", X"FA40", X"F95A", X"F8F4", X"F8C6", X"F780", X"F8A6", X"F625", X"F641", X"F683", X"F995", X"FCBC", X"FE8A", X"0295", X"FF5A", X"FE4A", X"FDC7", X"0088", X"005C", X"FCF6", X"FFF6", X"FBE9", X"FD74", X"FBC9", X"FC06", X"FC98", X"FBAC", X"FC35", X"FF6B", X"FE53", X"FCED", X"FCEB", X"FDD3", X"FBFD", X"FABD", X"FA9A", X"FB69", X"FD11", X"000F", X"013D", X"0270", X"FFAA", X"FF13", X"0095", X"FFAA", X"0010", X"FEB3", X"01A3", X"004B", X"FDA9", X"FEFB", X"FEDE", X"FDF3", X"0075", X"00CD", X"00D7", X"FF97", X"FFC6", X"004C", X"FFEA", X"FD7A", X"FEA3", X"000B", X"FEDF", X"008C", X"00FF", X"0405", X"0431", X"0295", X"0301", X"020D", X"0168", X"FEF7", X"0068", X"FF2D", X"032B", X"02B3", X"FDFE", X"FFDC", X"FF92", X"FE90", X"FF85", X"015A", X"012B", X"0094", X"015C", X"0201", X"01BE", X"FFBF", X"018D", X"0350", X"03AD", X"029E", X"056B", X"04F9", X"03F0", X"0266", X"00F7", X"0384", X"0146", X"FF4E", X"FDE6", X"0170", X"0264", X"004F", X"FCD2", X"FFF0", X"FF04", X"FDEF", X"FF99", X"018C", X"01EA", X"00A2", X"0071", X"FFF8", X"012B", X"0164", X"FFF4", X"0199", X"02B7", X"0301", X"02C8", X"0439", X"0341", X"0598", X"061A", X"07FA", X"FF4C", X"FF7F", X"00D2", X"022E", X"00FE", X"FFFB", X"FB98", X"FF88", X"FD3C", X"FBD7", X"FE50", X"FFB8", X"FE44", X"0216", X"011B", X"FFB9", X"FE71", X"011B", X"027F", X"03F5", X"0296", X"0210", X"015C", X"0352", X"02B5", X"03B9", X"0814", X"0950", X"01E9", X"0506", X"0012", X"04FA", X"0209", X"FE8E", X"FC06", X"FBA7", X"FCEB", X"FE19", X"FE7A", X"01A5", X"0194", X"016E", X"0286", X"0173", X"FE00", X"0352", X"02F7", X"0182", X"0214", X"0064", X"FE93", X"0050", X"0004", X"FE1E", X"0425", X"0BAD", X"07B1", X"02DB", X"01A9", X"006B", X"017F", X"FE8D", X"FCD2", X"FDFB", X"FF3E", X"FF67", X"015F", X"01C6", X"00D0", X"0396", X"03F3", X"00E6", X"FE5E", X"04BF", X"02DD", X"0062", X"FE23", X"FA48", X"F937", X"F966", X"F756", X"F435", X"F728", X"07EF", X"0373", X"0223", X"0235", X"0308", X"0723", X"FF86", X"00D1", X"FF8A", X"006F", X"02A5", X"0119", X"0133", X"0378", X"0409", X"0240", X"FF12", X"FDA4", X"0204", X"0320", X"FE62", X"FCDD", X"FB66", X"F8F7", X"F595", X"F2B2", X"EFCA", X"F0F5", X"FCE6", X"FCD9", X"FD3D", X"FF32", X"FF87", X"041A", X"00A2", X"05BC", X"0331", X"018E", X"03A4", X"0238", X"016D", X"035E", X"02FC", X"0064", X"FC97", X"FE72", X"FFE3", X"006B", X"013A", X"0090", X"00AF", X"FF6A", X"FDD1", X"F566", X"F077", X"F3FC", X"F99A", X"F932", X"FDE7", X"01A2", X"FFD9", X"00B9", X"02F9", X"08DB", X"03EF", X"01B8", X"02C3", X"021D", X"022B", X"023A", X"00C8", X"FDFD", X"FAB7", X"FD26", X"00E0", X"042D", X"03B4", X"0315", X"0418", X"041A", X"FECB", X"FB81", X"F8DB", X"F7CE", X"FCEB", X"F88D", X"FDA7", X"02AC", X"0124", X"FDD8", X"0200", X"059F", X"03E7", X"043A", X"0273", X"010C", X"0115", X"0125", X"FF0C", X"FB95", X"F904", X"FB73", X"0147", X"04F2", X"05CA", X"043B", X"05B2", X"0120", X"FFCC", X"FD10", X"FBDB", X"F946", X"FBB8", X"FE4E", X"FDB7", X"FF79", X"FEAD", X"FC43", X"FDEB", X"0269", X"024F", X"044B", X"0314", X"03CA", X"0054", X"FF26", X"FF29", X"FECE", X"FB38", X"FED8", X"042B", X"02B9", X"0656", X"0509", X"0366", X"014B", X"0090", X"FE5C", X"FC39", X"FC6B", X"FB7C", X"FDB6", X"FFED", X"000C", X"FE9E", X"FC09", X"FAE8", X"0135", X"02DE", X"048C", X"0282", X"025F", X"FF8B", X"FDF7", X"FF22", X"FE67", X"FFFB", X"02A1", X"06F5", X"04C0", X"0434", X"0525", X"015F", X"0170", X"FEFA", X"FE1A", X"FD4C", X"FC8E", X"FB73", X"FE7C", X"FEC7", X"003F", X"FF41", X"FF39", X"FA2A", X"00E5", X"011A", X"03C3", X"FFCA", X"FFD5", X"FEA9", X"FF17", X"FE4D", X"FFA1", X"00B6", X"0537", X"0296", X"0166", X"00BF", X"FFB0", X"0115", X"0095", X"FBE9", X"F81D", X"FC53", X"F856", X"F8D6", X"02EF", X"FE2E", X"0049", X"FCAB", X"FE61", X"FB3B", X"0216", X"007B", X"0229", X"FDE1", X"FD40", X"FC20", X"FC8E", X"FCA0", X"FCD5", X"003E", X"0114", X"FF68", X"FC52", X"FB81", X"FD19", X"FD97", X"FD73", X"F9BB", X"F72B", X"FBA7", X"FBD5", X"FDBE", X"FE88", X"FF8F", X"FEF2", X"FD03", X"FC51", X"F9A1", X"FD7B", X"FABC", X"FC99", X"F9F2", X"FC89", X"FBBB", X"F976", X"FC78", X"FA52", X"FBA2", X"FC24", X"FA6F", X"FB25", X"FB8F", X"FBB7", X"FBD1", X"FA04", X"F9DA", X"F8DD", X"FD56", X"020E", X"025F", X"FDDE", X"0013", X"FFBF", X"FE8E", X"F9C7", X"FCB6", X"FEC0", X"F91E", X"F80B", X"F93A", X"FB0D", X"FC4E", X"FC38", X"FAB8", X"FBB7", X"F984", X"F903", X"FAFF", X"FC92", X"FB17", X"FB49", X"FA42", X"F995", X"FBE0", X"FBFC", X"FDB1", X"058A", X"0441", X"FF28", X"FF37", X"FF83", X"002D", X"FA38", X"FEB1", X"FE52", X"F932", X"F8B6", X"FCDE", X"FF6E", X"0046", X"FF11", X"FE91", X"FE3D", X"FA1F", X"FA60", X"FC7E", X"FCB9", X"FBD2", X"FA23", X"FB60", X"FD8C", X"FDCE", X"FF3F", X"0244", X"06FF", X"037E", X"01F3", X"FF56", X"FF9D", X"FF48", X"FAFB", X"FEE7", X"0167", X"0078", X"FFB3", X"0016", X"007B", X"FECE", X"00BF", X"0031", X"FD24", X"FC08", X"FDB0", X"FE59", X"FD67", X"FAFF", X"FBE6", X"FD94", X"FF6E", X"004A", X"01A0", X"0401", X"048D", X"0310", X"00F1", X"007B", X"FF67", X"FF52", X"FF73", X"007F", X"0602", X"086F", X"0696", X"03C0", X"00A1", X"0095", X"0056", X"FD02", X"FD70", X"FC6A", X"FC8E", X"FCB1", X"FD15", X"FE0C", X"FC77", X"FE04", X"01A9", X"0486", X"0502", X"03F9", X"FF81", X"FC45", X"FDFB", X"FF91", X"0110", X"001B", X"FCF5", X"0435", X"07AA", X"093C", X"0644", X"0374", X"0178", X"FFB8", X"FDAE", X"FE12", X"FB99", X"FEBE", X"FDA9", X"FE0F", X"FF24", X"FF58", X"FF48", X"FF2A", X"036B", X"0505", X"0695", X"053C", X"03B3", X"FE30", X"FDE7", X"FFA8", X"009F", X"0026", X"FF37", X"FFDF", X"0398", X"0574", X"066F", X"03BE", X"03C2", X"063F", X"0448", X"061B", X"03DF", X"05DB", X"08AB", X"06DA", X"02E4", X"0393", X"03F1", X"051B", X"0335", X"0358", X"0319", X"01DB", X"FEB8", X"0031", X"0100", X"FFF3", X"009E", X"0154", X"FFC0", X"FF7B", X"FF3D", X"000F", X"FF7E", X"012A", X"0058", X"02F0", X"02FA", X"07E4", X"0495", X"062B", X"05D5", X"0766", X"0950", X"084E", X"033F", X"053E", X"0488", X"0323", X"03EC", X"02BE", X"0019", X"FE35", X"008D", X"FFE5"),
        (X"FF75", X"FF0D", X"0066", X"01C3", X"00AD", X"00C9", X"00D7", X"0154", X"FF63", X"FF84", X"004B", X"0052", X"FFB6", X"FF93", X"0068", X"014F", X"00D0", X"0075", X"FF84", X"0059", X"004E", X"FF69", X"00D6", X"0006", X"0003", X"FEDA", X"0041", X"0095", X"FF90", X"FEF4", X"0012", X"FF8B", X"FFA3", X"FF4F", X"FFF8", X"0035", X"FF8F", X"003A", X"FEA2", X"FF41", X"FF9F", X"FF65", X"0242", X"0225", X"FD91", X"FDEB", X"FD5F", X"FEBA", X"FE3C", X"FECE", X"FF01", X"0046", X"FE51", X"01C4", X"006E", X"002C", X"FF4E", X"000B", X"012C", X"FFEA", X"00B8", X"FEF2", X"0043", X"FCC3", X"FCFE", X"FE29", X"FB88", X"F8FC", X"F9F7", X"FD59", X"FEC3", X"FFB6", X"FFC7", X"FA72", X"FB81", X"FAFE", X"FD36", X"FCFA", X"FDE6", X"FCB8", X"FF7C", X"FE7F", X"0018", X"FF45", X"FFC1", X"00D5", X"0316", X"FE4B", X"FB3C", X"FE70", X"FD93", X"FB14", X"FB53", X"F79D", X"F6E4", X"F563", X"FA61", X"FC5B", X"FA03", X"FD64", X"FC35", X"F990", X"FC4F", X"F8D5", X"F9E3", X"FC74", X"FFAB", X"01BB", X"FFF1", X"0077", X"FBD5", X"FFB6", X"0078", X"0102", X"031B", X"01BC", X"00B2", X"FC19", X"FF42", X"FD56", X"FF05", X"FFCD", X"0053", X"003A", X"01A7", X"00F2", X"00EB", X"FEAF", X"FE7E", X"FB83", X"FB39", X"FD81", X"00E2", X"004E", X"00A6", X"FDB7", X"FD8F", X"011B", X"01DC", X"FEFC", X"FFB7", X"0047", X"027C", X"057B", X"FFAD", X"0152", X"0273", X"007C", X"001B", X"FE88", X"FF7E", X"020C", X"0315", X"032D", X"00A1", X"02C5", X"FED4", X"FD50", X"FCE0", X"FC93", X"FD5F", X"FBD5", X"FDDC", X"FD6A", X"FF6D", X"009E", X"008B", X"FD9E", X"00EF", X"FF07", X"FFCE", X"02FC", X"FCD8", X"FEC4", X"00C3", X"FF71", X"00F8", X"0119", X"0108", X"024F", X"02D6", X"0331", X"0059", X"0372", X"0261", X"02D2", X"0073", X"FFEF", X"0021", X"FEC0", X"FB61", X"FB30", X"FBFA", X"FFD8", X"FC90", X"0061", X"FEEC", X"FE4A", X"FFF2", X"0262", X"FF56", X"FF3C", X"017C", X"0104", X"01E7", X"01AF", X"022D", X"005C", X"004C", X"0301", X"0010", X"0433", X"03AC", X"00EE", X"0181", X"00C6", X"0275", X"001A", X"FC3E", X"FCCC", X"FCA9", X"FC94", X"FE24", X"FFBB", X"FE52", X"FE6C", X"0018", X"0415", X"01D6", X"019D", X"0202", X"0247", X"01C6", X"0183", X"0172", X"009D", X"0123", X"0001", X"020B", X"0195", X"0233", X"026B", X"028C", X"0378", X"0224", X"0098", X"00F4", X"FC8F", X"FBD7", X"FC80", X"FFFB", X"0287", X"0215", X"018B", X"0009", X"02A5", X"0233", X"0354", X"03DB", X"03D6", X"02DC", X"0191", X"0119", X"0125", X"009D", X"00B8", X"02C8", X"0543", X"02A6", X"0235", X"029E", X"02EF", X"0272", X"0181", X"FF91", X"FCC5", X"F956", X"F941", X"FBF2", X"0095", X"0044", X"02AF", X"02E8", X"0244", X"023A", X"055A", X"0467", X"03BF", X"0111", X"00D9", X"0224", X"009F", X"0003", X"01E4", X"0426", X"01F7", X"00EF", X"02F2", X"01CD", X"031B", X"0338", X"01BE", X"FFFC", X"FD71", X"F6FF", X"F6F2", X"F880", X"FF77", X"FF44", X"01DF", X"044F", X"04AC", X"0738", X"05C7", X"0560", X"03DF", X"02F5", X"02E5", X"005D", X"FE07", X"FD2D", X"007C", X"06A1", X"0408", X"01C7", X"028C", X"0479", X"0342", X"06AC", X"0892", X"0863", X"0257", X"FB8D", X"FC15", X"0002", X"0031", X"FFBA", X"0324", X"0449", X"0536", X"05E7", X"0497", X"028B", X"016C", X"008B", X"016A", X"FC84", X"FBB3", X"F97E", X"FFE7", X"0822", X"05A2", X"0388", X"03EF", X"0582", X"04FB", X"07F1", X"0BE7", X"0E87", X"08D3", X"0640", X"03D7", X"021D", X"00D3", X"FFAA", X"002B", X"0417", X"0245", X"06D2", X"0134", X"FE05", X"FED5", X"FED7", X"FC1D", X"FBA6", X"F8B2", X"FA62", X"0370", X"056B", X"07EA", X"05C0", X"029D", X"03E5", X"04BE", X"07AD", X"05DF", X"0582", X"03B0", X"FF0C", X"0194", X"01A1", X"FF18", X"FCB9", X"00C7", X"016E", X"0224", X"02FA", X"FF79", X"FBD4", X"FB51", X"FAF4", X"FA53", X"F993", X"FB87", X"FD5A", X"0411", X"0632", X"0616", X"031D", X"0222", X"00B7", X"FDDC", X"FE6F", X"FFB5", X"FD49", X"FCE3", X"FBE5", X"0038", X"FC2F", X"FD77", X"FE28", X"0358", X"FE9E", X"FF4D", X"0074", X"FC7A", X"FBF3", X"FB18", X"FAF8", X"FA7E", X"FA81", X"FB5C", X"FE1D", X"0382", X"056D", X"02C1", X"001E", X"FF02", X"FDEB", X"FBD6", X"FDAB", X"FA23", X"FAA5", X"F990", X"FAF5", X"FBA2", X"FB5D", X"FDBB", X"0128", X"0190", X"FF07", X"FE1B", X"FFAF", X"F993", X"FD77", X"FE0A", X"FFEF", X"FFF1", X"0032", X"FD3F", X"FF3E", X"0243", X"0214", X"006B", X"FD93", X"FC9D", X"FABF", X"FC0F", X"FA6E", X"F9B9", X"F952", X"FAE3", X"F786", X"F575", X"FACB", X"FE71", X"007A", X"02A4", X"FFC1", X"FE63", X"FDE1", X"F72F", X"F9B7", X"0080", X"0408", X"01EC", X"FEE1", X"FEC6", X"FF8A", X"01A8", X"FEFE", X"FD9E", X"FBA9", X"FCBC", X"FBAF", X"FB9A", X"FD3A", X"FC58", X"FA24", X"F8E9", X"F89F", X"F71C", X"FE28", X"0048", X"02BE", X"FFD9", X"03D6", X"FD16", X"F914", X"F66C", X"F8EA", X"FCB0", X"022E", X"02AF", X"0263", X"0018", X"FF40", X"FF3D", X"FE43", X"FB61", X"FC2E", X"FC75", X"FC66", X"FCFD", X"FD6C", X"FCBC", X"FA1C", X"F6A0", X"F47A", X"F716", X"0018", X"FE3C", X"FF80", X"01CC", X"0462", X"FC60", X"F86E", X"F908", X"F9E5", X"FD14", X"FEB0", X"FDFA", X"FE48", X"FBFD", X"FDCE", X"FD0F", X"FB4D", X"FBB8", X"FCC3", X"FCD5", X"FB92", X"FCD7", X"FCFF", X"FCC4", X"FB69", X"F840", X"F689", X"F9E5", X"FD8D", X"007E", X"0142", X"FD5F", X"FE02", X"FB9B", X"F905", X"FA51", X"FBEF", X"FD49", X"FCE4", X"FBBB", X"FD23", X"FADC", X"FBF5", X"FEEE", X"FE14", X"FCF9", X"FCCB", X"FE42", X"FE8A", X"FE29", X"FFE0", X"FC55", X"FB2D", X"F785", X"FA08", X"FF1A", X"FCFE", X"FFB1", X"019B", X"012F", X"FE34", X"FAFC", X"F9F3", X"FBA5", X"FCC1", X"FE9A", X"FCCB", X"FB6B", X"FD0C", X"FD47", X"FEB3", X"0016", X"0124", X"0257", X"00C0", X"FFEE", X"FE74", X"FFD8", X"00AF", X"FE53", X"FCE3", X"FA0F", X"FAB6", X"FF49", X"FC2E", X"FF7A", X"003F", X"024B", X"FF1B", X"FC5E", X"FB9C", X"FDA6", X"FFC6", X"FFA8", X"FF39", X"FCB2", X"FF50", X"FF55", X"007A", X"014D", X"048F", X"043D", X"0199", X"0195", X"01BF", X"005B", X"FFC6", X"FEEE", X"FE91", X"FC41", X"FAE9", X"FD11", X"FB2B", X"FFB5", X"FFF1", X"FF2A", X"FFA9", X"FCDA", X"FCAE", X"FC60", X"FDEE", X"009F", X"008B", X"0094", X"FEF7", X"0062", X"0165", X"038B", X"024B", X"0210", X"0408", X"02FC", X"0195", X"FF6C", X"FFF2", X"FFF6", X"00C2", X"0032", X"FEFA", X"FD48", X"FDDB", X"010B", X"00A8", X"0007", X"00C8", X"FE23", X"00AC", X"0242", X"02FE", X"0206", X"03AE", X"0278", X"0333", X"025B", X"0070", X"FE71", X"FDCF", X"FD06", X"FE98", X"FFD5", X"FF03", X"010F", X"025F", X"00EB", X"0237", X"00F3", X"FFB5", X"FC74", X"FE36", X"FECE", X"0011", X"0099", X"008E", X"FDC5", X"011D", X"06E8", X"058B", X"0491", X"0846", X"0807", X"04AC", X"02C5", X"04E3", X"00C7", X"01C0", X"0119", X"028D", X"0396", X"021E", X"0294", X"05BD", X"0491", X"FFB9", X"FFCD", X"FDB5", X"FE99", X"FE6D", X"FFAC", X"FFEA", X"0092", X"006C", X"FEF1", X"0178", X"03BA", X"05EB", X"0858", X"083E", X"07ED", X"090B", X"04AB", X"068A", X"068F", X"0A49", X"0613", X"0547", X"052E", X"04DF", X"0495", X"03BD", X"02A5", X"0305", X"0310", X"02EE", X"FFBC", X"0071", X"FF99", X"0053", X"FFC2", X"0010", X"005C", X"002B", X"01B2", X"02FB", X"02C8", X"035A", X"0268", X"00AA", X"FF94", X"00B4", X"0240", X"0646", X"0384", X"033A", X"042E", X"0501", X"041D", X"0363", X"0405", X"0354", X"0390", X"00A4", X"FFE4", X"0109", X"00BF"),
        (X"006D", X"FFDB", X"00CB", X"FFCD", X"FF2B", X"0096", X"0041", X"0116", X"FF44", X"0072", X"0115", X"001F", X"00EF", X"FFBB", X"0122", X"FFFF", X"0091", X"0052", X"0065", X"00B1", X"00B7", X"0054", X"002F", X"FFFD", X"FFBA", X"FED1", X"FF54", X"0007", X"FF3B", X"0040", X"005F", X"FFBD", X"0030", X"FF9B", X"FF12", X"0094", X"007C", X"0310", X"02E9", X"FDA1", X"FD24", X"FE8D", X"01DE", X"FF1B", X"0281", X"026D", X"01B2", X"FFEB", X"007C", X"003E", X"00AC", X"0086", X"0014", X"0111", X"FF85", X"FF13", X"00A3", X"0187", X"FF08", X"FE89", X"FF19", X"0005", X"00BA", X"FE5C", X"0144", X"0386", X"0597", X"04B8", X"0068", X"0335", X"0268", X"00A9", X"FF2B", X"00C6", X"0239", X"01EB", X"04BA", X"0718", X"0581", X"06F0", X"04A5", X"01EF", X"FFA9", X"0022", X"FF8B", X"FEA3", X"FE02", X"FD69", X"FDE4", X"FD65", X"FD9D", X"FF76", X"031F", X"04ED", X"05CD", X"053A", X"0479", X"050D", X"0257", X"012C", X"0380", X"0209", X"0217", X"0262", X"038C", X"02EB", X"0507", X"0167", X"027E", X"043C", X"0123", X"004A", X"014D", X"016F", X"FF70", X"FD50", X"0320", X"FF06", X"0084", X"01FC", X"04D9", X"07FB", X"0745", X"050C", X"0592", X"0204", X"00AE", X"FE40", X"027D", X"027B", X"00DC", X"01A8", X"006D", X"FEF9", X"FD04", X"FD35", X"FF24", X"01D3", X"FE0F", X"0172", X"0082", X"FF9E", X"FDDA", X"FE4A", X"032E", X"01DB", X"022A", X"04AA", X"081D", X"0944", X"08FF", X"064E", X"0208", X"01E2", X"0123", X"0110", X"02C8", X"031D", X"00FE", X"00EE", X"FF08", X"FF13", X"FCB9", X"FAFD", X"FC2D", X"02ED", X"FFD4", X"024B", X"FFCE", X"FFDB", X"FFB7", X"0067", X"007E", X"0406", X"031E", X"0469", X"0526", X"06EF", X"0603", X"0543", X"014A", X"FE24", X"FED8", X"FFCF", X"02A7", X"0094", X"FF63", X"FF75", X"FEAD", X"00A5", X"FE50", X"FDE6", X"FB5C", X"FE41", X"FE90", X"0058", X"00DC", X"0106", X"0387", X"0155", X"0608", X"0560", X"03FB", X"01FC", X"048F", X"0527", X"0366", X"0294", X"FEF3", X"FD15", X"FDDA", X"FFA8", X"FE75", X"FF19", X"FE4A", X"FD8A", X"FD33", X"00B8", X"0004", X"FCBC", X"FB5B", X"FB76", X"FF65", X"0074", X"FCBF", X"02BD", X"03E6", X"02F3", X"08C6", X"0480", X"026C", X"01B5", X"0296", X"028C", X"02C3", X"02F3", X"FEE9", X"FCB8", X"FDC9", X"FE91", X"FDC0", X"FEAA", X"FE2E", X"FD6C", X"FEF5", X"001B", X"FF4B", X"FE91", X"F85C", X"FAC4", X"FF09", X"FE2D", X"00B4", X"0300", X"05ED", X"041E", X"068F", X"029B", X"00AC", X"0114", X"00E5", X"033D", X"0325", X"0312", X"FF76", X"FD02", X"FD5B", X"FD68", X"0140", X"FE13", X"FE09", X"FDDD", X"FF12", X"01D1", X"00A9", X"FE82", X"F7A1", X"F820", X"FB7F", X"FF10", X"01C3", X"FFCA", X"04F1", X"0495", X"055C", X"034A", X"00A5", X"00EC", X"028F", X"03FC", X"04C2", X"015E", X"FDD8", X"FA70", X"FA8B", X"F9D0", X"FC6C", X"FD0D", X"FF90", X"FF0A", X"FEBF", X"FE92", X"00E5", X"FB5B", X"F603", X"F421", X"F885", X"001A", X"FF7C", X"00D9", X"02DA", X"054C", X"0706", X"045D", X"0101", X"FFFA", X"02C2", X"05BC", X"0586", X"01A3", X"FEEB", X"F844", X"F7F4", X"F879", X"FC33", X"FCFC", X"FE5A", X"0108", X"FF01", X"FE44", X"0061", X"FD33", X"F715", X"F727", X"FA12", X"FF2A", X"FF5D", X"0270", X"0438", X"05C4", X"01E4", X"FFFA", X"FEA0", X"00F4", X"04D7", X"0413", X"0473", X"030B", X"FE89", X"F9CB", X"F7F0", X"FA6B", X"0012", X"FF89", X"0146", X"0234", X"0229", X"FF92", X"0145", X"FEDA", X"0315", X"00FC", X"FD9E", X"0152", X"FFAA", X"007C", X"0337", X"01E7", X"FF9B", X"FEA7", X"FF15", X"00C4", X"0216", X"0436", X"04CC", X"02A2", X"FDA9", X"FD8D", X"FB2E", X"FDC6", X"02FB", X"048C", X"05FC", X"038A", X"0380", X"014A", X"FF0B", X"FEAD", X"055A", X"06E1", X"04FC", X"0178", X"FFC7", X"FEE8", X"0226", X"FF73", X"FCC8", X"FE48", X"FF1D", X"0340", X"02D2", X"0328", X"0363", X"03C8", X"0007", X"FF53", X"0105", X"0338", X"03F3", X"0615", X"0622", X"0616", X"034E", X"009F", X"FF63", X"FD05", X"FD49", X"07FF", X"061C", X"0111", X"FEEC", X"FEE7", X"FF15", X"00DC", X"FCB8", X"FD89", X"0076", X"0302", X"0292", X"0538", X"05DC", X"0510", X"02C9", X"028C", X"034D", X"041A", X"0353", X"0513", X"0405", X"071F", X"04AA", X"041F", X"FFED", X"FC97", X"FCD2", X"06A7", X"04C8", X"039A", X"00AE", X"FE6F", X"FDBB", X"FEE1", X"FCA0", X"FC0D", X"FBE6", X"0165", X"0649", X"07C4", X"076E", X"072A", X"07DE", X"05E4", X"0227", X"0190", X"0464", X"03CD", X"02C4", X"057D", X"062B", X"059E", X"0073", X"FB53", X"FEC2", X"08A5", X"059D", X"01F6", X"003F", X"FD53", X"00BE", X"FE7F", X"FD06", X"FB00", X"F9FD", X"FDB9", X"0282", X"0809", X"0867", X"0AC9", X"09C3", X"036B", X"FF79", X"FDC7", X"0150", X"0126", X"03B4", X"0716", X"050A", X"0328", X"FF66", X"FB2C", X"FDDB", X"06FD", X"02AB", X"009D", X"00AC", X"FF5B", X"018E", X"0086", X"FF8A", X"FDD4", X"FA61", X"F8FA", X"FB2B", X"01B8", X"04E8", X"0462", X"0354", X"FFF4", X"FB23", X"FB6B", X"003B", X"00E7", X"0363", X"06BE", X"0334", X"0385", X"FEDC", X"FED6", X"0083", X"00BD", X"01F1", X"FD09", X"FEC6", X"0086", X"FD82", X"FE5D", X"003F", X"FE02", X"FCC3", X"FB0D", X"FC15", X"FDFD", X"FF72", X"0186", X"011E", X"FE82", X"FBC8", X"FE17", X"FF7D", X"0190", X"03E8", X"0472", X"0437", X"0174", X"FE8C", X"FCDB", X"FDC2", X"FFBF", X"0103", X"FE33", X"01A4", X"FCFC", X"FE2B", X"FE9B", X"005C", X"FE05", X"FCBB", X"FE09", X"F97B", X"FA94", X"FD17", X"FEA6", X"00C4", X"FF20", X"FE11", X"FFB2", X"01C3", X"004C", X"02E5", X"03D7", X"038E", X"0222", X"FF0D", X"0090", X"009C", X"025A", X"0099", X"FF3D", X"FE6E", X"FFC1", X"00FA", X"010A", X"FFA1", X"FEEF", X"FBCD", X"FC6F", X"F9FC", X"FAB8", X"FC7F", X"FDD2", X"016A", X"0079", X"FF99", X"0129", X"0296", X"04BA", X"0585", X"0565", X"009C", X"FE46", X"FF10", X"03B9", X"04FA", X"01B2", X"0005", X"FF66", X"00DF", X"003E", X"022D", X"0490", X"0264", X"FFB0", X"0028", X"FDFE", X"FC40", X"F9DD", X"FC07", X"FF12", X"0055", X"0007", X"FF06", X"0219", X"0189", X"0463", X"055A", X"01F6", X"0169", X"0122", X"00B7", X"00CB", X"0531", X"FFED", X"FEE9", X"FF35", X"FE31", X"00EF", X"00FA", X"02D3", X"0384", X"FEE5", X"00DC", X"FEC1", X"FE63", X"FC1B", X"FD1D", X"FD98", X"FD3F", X"0119", X"03C7", X"02BD", X"01E4", X"0342", X"0365", X"0573", X"03B8", X"0473", X"060F", X"0205", X"0075", X"FE55", X"FE4D", X"0069", X"003A", X"FF91", X"FF21", X"01FD", X"0493", X"01F2", X"03B0", X"02AC", X"015E", X"00BE", X"00F0", X"0337", X"02AE", X"024B", X"03B1", X"026A", X"04C0", X"0268", X"03BB", X"02BE", X"03AD", X"03F9", X"0316", X"0080", X"001F", X"0097", X"FEFB", X"0105", X"000D", X"FF45", X"00C1", X"00A8", X"07AF", X"0647", X"06CF", X"093B", X"088E", X"0790", X"088B", X"0771", X"0603", X"0628", X"0820", X"0796", X"0531", X"03B8", X"03B1", X"01E6", X"0043", X"0011", X"01E1", X"00C9", X"0061", X"0123", X"0118", X"0136", X"0041", X"FFF1", X"001A", X"FD4C", X"FEB3", X"02BE", X"04D2", X"098E", X"0AA1", X"0657", X"04A1", X"055A", X"0272", X"0492", X"0598", X"0217", X"00EE", X"04F0", X"0326", X"0154", X"00ED", X"0281", X"0446", X"0460", X"0020", X"0067", X"FF8D", X"FF8D", X"FF2B", X"0003", X"0062", X"0067", X"01DA", X"01D2", X"035B", X"04B5", X"0473", X"02D8", X"04BF", X"0277", X"03BC", X"0576", X"0308", X"02DE", X"03B9", X"0274", X"029A", X"0430", X"0302", X"0420", X"02D9", X"037C", X"00B5", X"00B4", X"FFCE", X"0058"),
        (X"001B", X"FFE1", X"0101", X"FF7C", X"001F", X"0002", X"0110", X"FFB2", X"FFDE", X"00B3", X"FFCA", X"004D", X"FE2F", X"FEB6", X"0075", X"01B4", X"001F", X"FF4E", X"FF89", X"FFC8", X"0051", X"FFA8", X"018C", X"FFC6", X"FF17", X"0065", X"FF0A", X"FF4C", X"FF6F", X"0171", X"FE9F", X"007E", X"FF3A", X"FFB8", X"008A", X"FE59", X"FEC2", X"FD19", X"FE46", X"FFD8", X"00EE", X"0046", X"FD07", X"FDB3", X"0220", X"0147", X"FCBF", X"FD1D", X"FD10", X"FCB6", X"FBA9", X"FF00", X"FF4C", X"FF71", X"FEEC", X"FFF0", X"0060", X"008E", X"FE29", X"01F1", X"0073", X"FF5F", X"FD92", X"FEBE", X"FEF8", X"FD48", X"FEFD", X"FEB6", X"FA8F", X"F865", X"F9CF", X"F901", X"F9E0", X"FB44", X"FE46", X"FC9E", X"FD94", X"FBEF", X"FBAD", X"FD86", X"FE2C", X"00AA", X"0039", X"005D", X"FF07", X"FF65", X"FFA6", X"0027", X"0001", X"FDC7", X"FC8F", X"FD77", X"FFC2", X"FF12", X"009A", X"0332", X"0034", X"00DA", X"FE3C", X"FDA3", X"FF2E", X"FFBB", X"01C6", X"FF3D", X"FE6D", X"FD14", X"FC63", X"FD61", X"FA65", X"FDA3", X"FF18", X"0083", X"FF1E", X"0105", X"FF82", X"008F", X"FDED", X"FD5F", X"0112", X"FD73", X"007D", X"01C2", X"0254", X"03EA", X"0123", X"0071", X"0018", X"018F", X"0223", X"0249", X"0319", X"FF44", X"FE1C", X"FDAA", X"FE43", X"FB15", X"FF8D", X"FF81", X"02AA", X"0008", X"0070", X"019A", X"FECA", X"03A2", X"FF2C", X"FCA9", X"FC25", X"FD86", X"FD2A", X"FE3E", X"006F", X"01FE", X"FF70", X"0217", X"0165", X"00D5", X"037A", X"0705", X"0544", X"0212", X"018E", X"FFBB", X"FE85", X"FB4F", X"FD1B", X"FF61", X"00D6", X"FE18", X"FFB8", X"FEEE", X"0139", X"FF6E", X"FECB", X"FC32", X"F9B9", X"F918", X"FA53", X"FC2A", X"FC14", X"FDE2", X"00A2", X"0489", X"03E7", X"0552", X"05FA", X"065E", X"05CE", X"02A7", X"032A", X"008B", X"FDFA", X"FDD2", X"FD94", X"FEC8", X"FF27", X"FFDF", X"003F", X"FD7B", X"FD4F", X"FCEA", X"FD17", X"F99A", X"FBE9", X"F915", X"FB41", X"F927", X"FBBB", X"FF8F", X"02D8", X"05D8", X"0669", X"07BE", X"0676", X"036B", X"02A2", X"00DF", X"0261", X"0060", X"0043", X"FEAC", X"FF9F", X"0259", X"FE8B", X"FF73", X"011B", X"FAFA", X"FBB9", X"F965", X"FC6B", X"FD29", X"FD2E", X"FB2F", X"FD3E", X"FD9F", X"FFFA", X"FD31", X"0060", X"01CE", X"035C", X"05C4", X"0717", X"0476", X"0365", X"021D", X"0033", X"FF8E", X"FF19", X"0018", X"0387", X"0385", X"023A", X"01AD", X"FF99", X"FA8B", X"F9BC", X"FAF8", X"F99B", X"FC0A", X"FD96", X"FE86", X"FE28", X"FEF6", X"FF2E", X"FD87", X"FF9F", X"002E", X"01B1", X"0139", X"027B", X"02D6", X"01D1", X"022C", X"FF75", X"FE13", X"FF33", X"0221", X"06AB", X"0581", X"0656", X"FFF2", X"FE6A", X"FAC5", X"FA20", X"FB4E", X"FAC8", X"FDAE", X"FF6C", X"FD9D", X"FF6E", X"FDD0", X"FDC3", X"FEBF", X"009E", X"00CB", X"0133", X"FF4D", X"FF20", X"0221", X"0258", X"0075", X"FF2A", X"FE90", X"FEFC", X"03FD", X"0753", X"06E8", X"07DD", X"FFC8", X"FEFD", X"FBAF", X"F8BE", X"FB29", X"FAA4", X"FE7C", X"FF6D", X"FE87", X"0055", X"FE9B", X"FE39", X"FF56", X"0071", X"0440", X"022F", X"FF7A", X"FE8F", X"0097", X"FFE0", X"0169", X"0333", X"01A1", X"01AE", X"03BF", X"05E6", X"068C", X"06E5", X"FF3B", X"FD5C", X"FA32", X"F755", X"F99B", X"FAD1", X"FC90", X"FFB2", X"FDC9", X"FCF4", X"FEF4", X"FF2A", X"0284", X"04B6", X"0796", X"0576", X"FFB2", X"FD16", X"00F3", X"003F", X"01C4", X"02F2", X"0138", X"01AF", X"01D0", X"FF6E", X"FEFF", X"03A3", X"FE4F", X"0057", X"FD77", X"F9CC", X"FA12", X"FDB3", X"FFFD", X"FF06", X"FCD5", X"FDE0", X"005E", X"0151", X"030B", X"06E2", X"0A16", X"0236", X"FC62", X"FDE6", X"FF88", X"007B", X"FFCC", X"FF70", X"FF87", X"FEEB", X"FED1", X"FC50", X"FDD2", X"033D", X"03D5", X"FE3F", X"FDF5", X"F999", X"FE14", X"FDEC", X"FE59", X"FDA2", X"FDDF", X"FEC1", X"02F2", X"0491", X"05CA", X"05EE", X"046F", X"FFBC", X"FCE1", X"FE51", X"FEFB", X"FD48", X"FB7C", X"FE6D", X"FF04", X"FCEA", X"FCB8", X"0130", X"FFC0", X"05B0", X"02F2", X"0010", X"0191", X"FA76", X"FC9F", X"012E", X"FFE9", X"FBEE", X"FF23", X"FFD0", X"0567", X"0867", X"0829", X"0543", X"FEB6", X"F9B6", X"FB2D", X"FE25", X"FD5C", X"FCED", X"FE03", X"FCD4", X"FE06", X"FBA8", X"FE58", X"01A3", X"007E", X"073F", X"018B", X"FE87", X"0058", X"FEAD", X"FE41", X"018D", X"02AB", X"FE17", X"FEE4", X"034D", X"07B4", X"0A02", X"095B", X"03DA", X"FB6A", X"F8B8", X"F9B7", X"FC7D", X"FDBB", X"FE66", X"FF23", X"FF67", X"FCA9", X"FF02", X"0093", X"012A", X"01EF", X"0906", X"0176", X"005C", X"FFC6", X"FF29", X"0017", X"03DB", X"0263", X"0213", X"055D", X"0793", X"0A36", X"0A46", X"0771", X"008C", X"FA53", X"F7DD", X"FA6E", X"FD47", X"FEEB", X"FE4C", X"FFF7", X"001F", X"FEB7", X"FE25", X"003C", X"FECD", X"FF6E", X"03A8", X"02F9", X"FDE7", X"FFB8", X"FE7F", X"FFE0", X"0529", X"03C5", X"067E", X"075D", X"09F9", X"0B8A", X"09BA", X"03A2", X"FADB", X"F807", X"FA9F", X"FD0E", X"FE9E", X"FF3D", X"0044", X"020A", X"0085", X"011D", X"01D3", X"01E8", X"FF32", X"002D", X"FF63", X"FF28", X"FFB7", X"FDBB", X"FE53", X"049A", X"0619", X"07FE", X"068C", X"065A", X"09C4", X"083E", X"042F", X"FE40", X"FA0B", X"FB3B", X"FAC9", X"FAAD", X"FCB5", X"0198", X"03BD", X"040F", X"032A", X"0383", X"053D", X"0481", X"0296", X"0320", X"024F", X"FD3E", X"FEE5", X"0095", X"0105", X"050C", X"09BA", X"09A5", X"080A", X"06FD", X"0632", X"0466", X"0081", X"FC90", X"F97B", X"F8B5", X"F8CF", X"FBC4", X"FD65", X"FF80", X"006A", X"02C4", X"0451", X"0408", X"0808", X"0615", X"060F", X"07DA", X"008B", X"FEF9", X"005F", X"00FB", X"0323", X"066E", X"09B1", X"06B4", X"06FD", X"0490", X"0153", X"00D7", X"FF2E", X"FCB4", X"FD69", X"FDB5", X"FBA7", X"FBA5", X"FC69", X"FE65", X"FFF0", X"002D", X"01DB", X"0342", X"07A8", X"071C", X"0527", X"0491", X"0168", X"FF6E", X"FF81", X"FEFB", X"026D", X"0793", X"05FE", X"035C", X"046A", X"017E", X"0007", X"01E6", X"0221", X"03D7", X"038F", X"032A", X"FFB0", X"FF8E", X"FE9A", X"FF24", X"002F", X"0069", X"0338", X"0302", X"06BD", X"0808", X"048C", X"FFDC", X"FFBE", X"0021", X"FF86", X"FEDD", X"03CC", X"07C7", X"047D", X"0199", X"FE55", X"FDF8", X"033B", X"023D", X"058E", X"0578", X"0389", X"0374", X"0284", X"0095", X"FF1E", X"FD40", X"01FA", X"00F0", X"01B1", X"0573", X"0640", X"08A8", X"0525", X"007E", X"FE52", X"FED0", X"012B", X"00C9", X"0104", X"02C4", X"FFC7", X"FCCD", X"FF36", X"FFD8", X"0139", X"00DE", X"0292", X"FFFF", X"FF8B", X"0068", X"0077", X"0300", X"0106", X"01F4", X"02B1", X"045E", X"0463", X"03F3", X"0696", X"07DE", X"02AA", X"0033", X"FDFB", X"FFB1", X"009D", X"0031", X"021F", X"FC98", X"FE12", X"00B7", X"0070", X"033D", X"00ED", X"0064", X"04A0", X"00E5", X"0167", X"0036", X"FF89", X"0176", X"0310", X"0270", X"039F", X"0563", X"057D", X"0697", X"01DE", X"0376", X"02D7", X"0325", X"0146", X"0179", X"FFDF", X"012D", X"FF09", X"0138", X"04D0", X"031E", X"025F", X"0206", X"03BC", X"0342", X"04DB", X"0447", X"03A6", X"045E", X"064A", X"0182", X"01C6", X"0143", X"0136", X"FEA4", X"0261", X"023A", X"FFE9", X"FF45", X"00AC", X"003A", X"FF69", X"FF40", X"008E", X"FF06", X"002C", X"FFA1", X"FF1F", X"FE2E", X"00AA", X"009E", X"0073", X"01F8", X"00E6", X"0138", X"FFE7", X"F94E", X"0070", X"FE17", X"FAB9", X"FA4C", X"FBD8", X"FC8F", X"FE3E", X"FE7B", X"FFE8", X"FB75", X"FF4E", X"0017", X"000E", X"FF4C"),
        (X"0069", X"FFEF", X"FE8D", X"010A", X"005B", X"FF03", X"FEDE", X"0102", X"FFE4", X"00BF", X"FF54", X"007B", X"0244", X"01AB", X"0103", X"FF91", X"00F0", X"FF27", X"00FA", X"0135", X"FF95", X"0083", X"00BA", X"FF4F", X"FEDF", X"FF92", X"FF5E", X"FFE5", X"FFB4", X"FEAB", X"00DD", X"FF26", X"FFC8", X"003D", X"0492", X"0565", X"044A", X"0424", X"0422", X"05D4", X"0592", X"05B8", X"047A", X"04DC", X"03EE", X"0546", X"02C8", X"033A", X"03D8", X"032F", X"03D5", X"02AC", X"01BD", X"FF3B", X"0035", X"00F7", X"FFD4", X"FF86", X"FFD5", X"0156", X"01FE", X"00B9", X"05EC", X"074F", X"09F0", X"0A38", X"0BA3", X"0DE7", X"0DAD", X"0E11", X"0F09", X"0B27", X"0863", X"05E7", X"0271", X"0046", X"0262", X"0432", X"0516", X"04A3", X"0374", X"01C8", X"00DB", X"FFE2", X"00C8", X"0015", X"FF96", X"03F8", X"0049", X"01F4", X"050F", X"0992", X"06AF", X"0A58", X"07A3", X"095F", X"06CC", X"0A15", X"07BA", X"0726", X"0614", X"0313", X"FB46", X"FD80", X"FC49", X"FC27", X"FC3B", X"FD22", X"FDF8", X"0413", X"0362", X"FF5C", X"FFED", X"FFD6", X"FECA", X"FD39", X"FFF7", X"FF4A", X"FF72", X"008B", X"FE20", X"FE2B", X"FE88", X"FF50", X"02E8", X"02EC", X"01F9", X"0075", X"FDFF", X"FDC9", X"FB52", X"FBC8", X"FC7D", X"FCA4", X"0070", X"FE46", X"FAC8", X"F793", X"FB06", X"02AA", X"005D", X"FEEF", X"0148", X"0198", X"01D0", X"FCF9", X"FD23", X"FCA2", X"FBD5", X"FC11", X"FC3D", X"FCAE", X"013D", X"02F8", X"02AA", X"04AF", X"027E", X"0102", X"0205", X"02BD", X"011F", X"02F2", X"0233", X"00D1", X"FE59", X"F9A9", X"FD13", X"005D", X"001C", X"FD0D", X"FF41", X"0163", X"042F", X"FE25", X"FE1C", X"FD6D", X"FAD3", X"FA62", X"FA15", X"FA9F", X"004F", X"02DD", X"0363", X"01D8", X"01A6", X"FF0A", X"00E0", X"0287", X"0237", X"02B2", X"030D", X"0012", X"FCF1", X"F901", X"FA15", X"FFC3", X"FFC0", X"FC10", X"FF69", X"FD67", X"FEF6", X"FDBF", X"FE4F", X"FE15", X"F988", X"FA12", X"FBA4", X"FBCD", X"FF3A", X"020F", X"039C", X"FED8", X"FEA8", X"FE6B", X"0058", X"FE75", X"FD0C", X"0114", X"00AB", X"FD63", X"FA14", X"F7C4", X"FCB6", X"0100", X"0228", X"FF55", X"0104", X"FE02", X"FF22", X"FE0C", X"FC0E", X"FBE7", X"FA98", X"FD77", X"FC00", X"FDFD", X"FE9E", X"02C9", X"0374", X"01F1", X"0015", X"FF53", X"FD6B", X"FE4C", X"FE0C", X"FD51", X"FC0C", X"FD28", X"F58E", X"F0F9", X"F76E", X"FBA1", X"FFA1", X"FD00", X"01EF", X"FEE7", X"FD7A", X"FE1D", X"FCAF", X"FCCF", X"FCC9", X"FD73", X"FCFC", X"FCA8", X"00A0", X"067C", X"0789", X"03B2", X"010C", X"0083", X"0091", X"0009", X"FCF2", X"FB04", X"F92D", X"F8CC", X"F5B7", X"F175", X"F66C", X"FBDA", X"009C", X"0064", X"FF2A", X"FE41", X"FBC6", X"FEF7", X"FC0F", X"FB3A", X"FE5B", X"FD62", X"FCFA", X"FB89", X"FDD1", X"02FE", X"0583", X"0377", X"FF55", X"014D", X"016A", X"00B3", X"FE1E", X"FC69", X"F9F5", X"F9BE", X"F858", X"F084", X"F6A6", X"FCD0", X"FFC1", X"02BC", X"FD34", X"0182", X"FBE1", X"FC9C", X"FDA2", X"FABB", X"FD0A", X"F9F1", X"FAEB", X"F933", X"F903", X"FDAF", X"0104", X"FF0C", X"FB47", X"FC4C", X"FF04", X"01CB", X"FEDD", X"0015", X"FE44", X"FF88", X"FCAD", X"F5EF", X"F560", X"FE04", X"FFD7", X"FDF9", X"FC29", X"FF9D", X"FC9A", X"FB5A", X"FD49", X"FC55", X"F9FC", X"F951", X"F7E1", X"F98D", X"FADD", X"FA98", X"FDF2", X"FED0", X"FB54", X"FD8E", X"FF1B", X"0253", X"0246", X"00FC", X"0011", X"04FB", X"05C8", X"0038", X"FC48", X"010B", X"014D", X"FE09", X"FF24", X"FF07", X"FE51", X"FC69", X"FD40", X"FBF9", X"FA86", X"F989", X"F898", X"F951", X"FBCD", X"FAEB", X"000E", X"FDEF", X"FD4B", X"FD61", X"007D", X"0119", X"002C", X"FE89", X"FF16", X"04B9", X"07A1", X"04EC", X"0508", X"02FD", X"FEBA", X"FD28", X"FE4D", X"0043", X"023C", X"0068", X"026C", X"02D9", X"FF7A", X"FC90", X"FAAF", X"FA70", X"F9B1", X"FD9E", X"0039", X"FFBB", X"FC50", X"F9BD", X"FD48", X"004E", X"00C7", X"FF64", X"FE0E", X"0176", X"0315", X"0677", X"07A6", X"027E", X"010C", X"FF7A", X"FFF0", X"FE81", X"0632", X"0822", X"05FF", X"04D3", X"0308", X"FF18", X"FD72", X"FA48", X"F9DE", X"FBDC", X"FF4A", X"FE56", X"FB11", X"F895", X"FE78", X"025E", X"0168", X"FEC9", X"FBED", X"FD67", X"030F", X"0873", X"021D", X"03CA", X"005D", X"FE8C", X"FF68", X"0118", X"0629", X"093C", X"0852", X"0681", X"02E4", X"02AC", X"029C", X"000D", X"FB77", X"FBA7", X"00F1", X"FC77", X"FB92", X"FBB3", X"0105", X"0440", X"0268", X"0174", X"0066", X"FE2E", X"0096", X"09C6", X"04F7", X"0334", X"FEEE", X"FC0C", X"FEDB", X"00D9", X"0676", X"0597", X"03B4", X"055E", X"05F7", X"0760", X"096A", X"0592", X"FF82", X"FEC2", X"0251", X"FE46", X"FC1D", X"FE1A", X"0198", X"020B", X"0271", X"007C", X"007D", X"FDFA", X"0030", X"0A14", X"04D2", X"053E", X"FEF3", X"FF4E", X"FDC0", X"FF00", X"0342", X"0142", X"03F2", X"03F1", X"05BF", X"0888", X"08EF", X"04D1", X"0372", X"0149", X"0455", X"01DB", X"FFEC", X"0216", X"046D", X"01F5", X"00A9", X"00BD", X"006A", X"0062", X"03E2", X"0894", X"0020", X"033E", X"0074", X"000B", X"FCCD", X"FBAD", X"FE20", X"FF15", X"0187", X"04A8", X"053A", X"0667", X"06C7", X"073C", X"07FA", X"07C2", X"0627", X"0353", X"034D", X"02E1", X"038C", X"0077", X"00AC", X"00FE", X"008D", X"0060", X"04F2", X"06E8", X"03D1", X"011B", X"00DE", X"011A", X"FD93", X"FC35", X"FE59", X"FED9", X"033B", X"0193", X"00C5", X"0257", X"03D8", X"05E1", X"0598", X"03D5", X"060E", X"02E6", X"0188", X"02A9", X"0332", X"0141", X"019B", X"018E", X"00D5", X"0045", X"0440", X"06BC", X"03CF", X"FFA5", X"000F", X"FE6F", X"FCAF", X"FD49", X"FC94", X"0135", X"0137", X"01DC", X"0079", X"0160", X"046B", X"026F", X"0423", X"0180", X"029A", X"015D", X"0169", X"0295", X"03F2", X"0489", X"0318", X"0349", X"03C4", X"0470", X"05E8", X"071F", X"0464", X"0024", X"FF06", X"0022", X"FDC2", X"FFEB", X"FB86", X"026E", X"01BF", X"021F", X"01E9", X"02E9", X"0288", X"009D", X"0011", X"FEFE", X"00D9", X"0010", X"0283", X"0316", X"03C8", X"028F", X"0126", X"0512", X"046B", X"04D6", X"04C3", X"05DA", X"00E6", X"00BF", X"FF7F", X"001E", X"FC8A", X"F898", X"F9DA", X"0101", X"FFCB", X"FFA7", X"010C", X"015E", X"00B8", X"00F5", X"0014", X"0014", X"FF78", X"FF57", X"01B0", X"037D", X"0443", X"01FE", X"02BC", X"04C5", X"05E6", X"0279", X"0376", X"052B", X"0173", X"00B4", X"001A", X"FFA9", X"FD89", X"F7A6", X"F674", X"F92A", X"F9E1", X"F9B7", X"FDA5", X"FF45", X"FBCC", X"FA92", X"FD74", X"FCFA", X"FD13", X"FE76", X"FE74", X"FFDB", X"FF9F", X"FC2C", X"FD72", X"00B0", X"015D", X"0005", X"040D", X"04CB", X"026B", X"FE54", X"FF1D", X"FFF1", X"00BF", X"FB99", X"FAA6", X"F4DA", X"F2DE", X"F392", X"F542", X"F3BE", X"EECE", X"F176", X"F12A", X"F214", X"F1AC", X"EEF4", X"EDE4", X"EF11", X"F24D", X"F6E4", X"F986", X"FB7A", X"FB3E", X"F9F3", X"FC91", X"0261", X"0334", X"00E6", X"FFD7", X"0094", X"0056", X"0003", X"FCF4", X"FD0E", X"FBA2", X"FABC", X"F84C", X"F91B", X"F80A", X"F9A6", X"FC0C", X"F6E0", X"F756", X"F914", X"F80F", X"F706", X"F9C7", X"0018", X"FE98", X"FC35", X"FC6C", X"FD9A", X"0389", X"FFCC", X"FEEF", X"00C7", X"FE15", X"01E1", X"00CB", X"0013", X"0015", X"FF46", X"FFBB", X"FFD3", X"FF94", X"FEDD", X"FD1C", X"FD9E", X"FEA9", X"FD92", X"FB90", X"FC78", X"FACE", X"FF2A", X"0032", X"FC30", X"FF1E", X"FD0C", X"FC17", X"FC09", X"FEBE", X"018E", X"00E2", X"00AA"),
        (X"FF25", X"FF1F", X"FF42", X"FEE2", X"FF6D", X"00B8", X"0045", X"FF7A", X"000C", X"0125", X"0004", X"007D", X"007F", X"016F", X"FF2A", X"000D", X"FFE4", X"00D1", X"0035", X"FFC9", X"FF3F", X"000D", X"00F6", X"00B9", X"007F", X"0096", X"FF2C", X"FFB0", X"00D9", X"003A", X"008C", X"FFFB", X"FFD6", X"0124", X"0207", X"033A", X"02D0", X"0250", X"02A5", X"0413", X"06CB", X"03B4", X"00CD", X"011C", X"FEF0", X"02BE", X"04C1", X"03DA", X"0435", X"0443", X"02C0", X"014F", X"00D7", X"0089", X"FF4D", X"FFB9", X"FF37", X"FF2A", X"00E8", X"014C", X"FFAF", X"007D", X"03E3", X"05D1", X"0322", X"00A8", X"0587", X"01FD", X"01AE", X"0161", X"0026", X"FF27", X"FEC0", X"000D", X"0185", X"0558", X"05C7", X"05AA", X"08BE", X"054E", X"0079", X"FCBC", X"FEC7", X"FFBD", X"0093", X"0025", X"FEC4", X"0094", X"02CC", X"FFA4", X"0120", X"01BB", X"FFF1", X"FED3", X"FCB2", X"FC3E", X"F999", X"FBF9", X"FB23", X"F980", X"F93C", X"FC52", X"FC94", X"FEAD", X"FE47", X"0214", X"0808", X"0A46", X"0679", X"02A9", X"03A3", X"FEC6", X"000A", X"0152", X"FEEA", X"FD75", X"0067", X"FDA3", X"FAEB", X"FD86", X"FE5A", X"FDDB", X"FD91", X"FEF4", X"FEC9", X"FDEF", X"FDAC", X"FE4A", X"FCD7", X"FD90", X"FDEF", X"00DF", X"006F", X"041A", X"0445", X"0AEF", X"09DD", X"0358", X"033F", X"0388", X"00B6", X"00FD", X"FF1D", X"FDCE", X"FF73", X"FA3E", X"FCD5", X"FC41", X"FF36", X"FE20", X"FF7C", X"FEE5", X"0123", X"020D", X"00CD", X"FE50", X"FC7D", X"FEDA", X"FFA7", X"FFA4", X"FF7E", X"0145", X"01AF", X"0482", X"07E5", X"0684", X"04A2", X"03A6", X"FFC3", X"FEAB", X"FD12", X"F97D", X"FBDF", X"F9C8", X"FDFC", X"FF8B", X"FE4E", X"FD4D", X"FDAC", X"FEF3", X"0014", X"006D", X"00F9", X"FFC7", X"FEBE", X"FDC6", X"FD2C", X"FEDF", X"FF45", X"FF3A", X"0174", X"0552", X"0705", X"086E", X"01BC", X"021C", X"0051", X"FCB0", X"FC47", X"F864", X"F9E7", X"FB55", X"FC8F", X"FD91", X"FE04", X"FC17", X"FBB7", X"FD20", X"FDEB", X"FCC8", X"FDB5", X"FED4", X"FE0E", X"FCFB", X"FDAE", X"FCF5", X"FD8E", X"FF57", X"FFFE", X"0572", X"0B3F", X"0BE3", X"0248", X"024C", X"0018", X"FE17", X"FB0B", X"FAC1", X"FBED", X"FDA9", X"FE25", X"FD2A", X"FC27", X"FB62", X"FBFC", X"FB76", X"FCFA", X"FFF7", X"0057", X"FD43", X"FE63", X"FC38", X"FCEF", X"FD4C", X"FF01", X"00E9", X"FD8D", X"04D0", X"0EE6", X"0C11", X"03A3", X"0038", X"0055", X"FE68", X"FBF2", X"FBF0", X"FE57", X"FDEC", X"008C", X"FF49", X"00A5", X"FEBB", X"0167", X"046B", X"0644", X"0C0E", X"08D3", X"00AB", X"FAA8", X"FBC0", X"FEA2", X"FFB0", X"0061", X"000F", X"0032", X"0296", X"0CB1", X"073E", X"036E", X"FF19", X"FEE6", X"0040", X"FACD", X"FD97", X"01C2", X"0304", X"05A9", X"07B4", X"071D", X"0907", X"0B8B", X"0FD4", X"11B6", X"11A5", X"0CB2", X"018E", X"FA89", X"FCCC", X"FED2", X"0063", X"0107", X"010A", X"02D5", X"0120", X"0554", X"FF43", X"FF4D", X"FE97", X"FFC6", X"FD9C", X"F9F9", X"FD6F", X"0673", X"0A1B", X"0ADD", X"0BDC", X"0FD7", X"1139", X"0FD0", X"0D70", X"0DBF", X"0D85", X"0859", X"001B", X"FC31", X"FDB1", X"FF02", X"FF44", X"00DD", X"0302", X"0437", X"0271", X"FFD8", X"FC3A", X"021C", X"019E", X"0015", X"FDF1", X"FCD2", X"009A", X"09D9", X"1012", X"0FDF", X"10A9", X"0F85", X"0E37", X"0AFA", X"05CE", X"0237", X"050F", X"05B8", X"0154", X"FECD", X"FE86", X"FFFE", X"01B6", X"03CC", X"04B5", X"0409", X"0441", X"FF0A", X"F9D3", X"F8C1", X"01A0", X"0022", X"FF4D", X"FDF8", X"03FE", X"0BC1", X"0FDE", X"0D62", X"0DA8", X"067C", X"04F7", X"02E8", X"FFA6", X"FF14", X"0031", X"04DC", X"0243", X"FF74", X"00BC", X"FFCC", X"014D", X"024A", X"0055", X"0523", X"01A6", X"FECB", X"F949", X"F9B2", X"FED5", X"021B", X"001E", X"FE93", X"047A", X"045D", X"09B4", X"0547", X"0198", X"0086", X"FDB7", X"FDA9", X"FE92", X"FDC2", X"FDF7", X"0010", X"00A4", X"FF07", X"FE90", X"006C", X"FE42", X"00A6", X"FD83", X"012B", X"011F", X"0048", X"F8D8", X"F775", X"FDF5", X"010D", X"FEA1", X"000F", X"0042", X"FE6E", X"000A", X"FDFC", X"FE03", X"FE9B", X"FE47", X"0052", X"FD93", X"FE46", X"FEE5", X"FF71", X"FE05", X"00EA", X"FFCA", X"014C", X"FFCE", X"00C9", X"FEC4", X"01CF", X"00B5", X"FB4E", X"FB81", X"FA3E", X"FDAA", X"FF36", X"FDF6", X"FCFF", X"FC51", X"FC30", X"FDC2", X"FC8F", X"FC53", X"FE5E", X"FE7A", X"FF7E", X"FE9B", X"FBC4", X"FE51", X"FEB1", X"FEFE", X"FF97", X"0081", X"0019", X"FD23", X"FFA2", X"FF9D", X"013D", X"01B5", X"FD49", X"F95E", X"F68D", X"FD2A", X"FFE1", X"FDFE", X"FC44", X"FC6F", X"F97A", X"FB4F", X"FCE3", X"FD63", X"00D4", X"FF3A", X"00B0", X"0024", X"FD5B", X"FF01", X"FFFE", X"0002", X"FFA5", X"FFCD", X"FEA8", X"FE1D", X"028D", X"01D3", X"02DC", X"01D9", X"FE20", X"FC36", X"FA6A", X"FD68", X"FF57", X"FEF5", X"FBD8", X"F822", X"F8F5", X"F9A1", X"FB8B", X"FD52", X"FF3B", X"012F", X"033D", X"01E7", X"FF65", X"FE90", X"0051", X"FE09", X"FF5B", X"FE20", X"FF64", X"FE6D", X"00B9", X"001C", X"0119", X"FFA2", X"FFB2", X"FC10", X"FAA1", X"FD13", X"006A", X"00EC", X"FF32", X"F9C8", X"FB35", X"FA39", X"FC58", X"FE3D", X"FFAF", X"00AD", X"0097", X"0117", X"00AE", X"FE92", X"FDC1", X"FDBA", X"FDA6", X"FE70", X"FFFD", X"FF35", X"0004", X"0143", X"FF23", X"FF4F", X"FD8A", X"FC5B", X"F9C6", X"FE2A", X"0023", X"0209", X"FCD4", X"F95B", X"FB46", X"FC1B", X"FD8B", X"FE70", X"011A", X"FEC4", X"00FB", X"FF03", X"018D", X"FFD4", X"FFA2", X"FFDC", X"FFF8", X"00E3", X"FE2E", X"0160", X"FEC3", X"00DA", X"0156", X"016D", X"FF29", X"FE5E", X"FB9C", X"0230", X"FFE3", X"FFB2", X"FB27", X"F999", X"FC84", X"FD52", X"FEB8", X"FF4F", X"FEC4", X"FFE2", X"0009", X"00A2", X"FEC8", X"0140", X"00FA", X"016D", X"0120", X"FF26", X"FFBC", X"FD48", X"01CC", X"0013", X"000D", X"FFF5", X"FDFF", X"FEAD", X"FCF7", X"FF6A", X"FFE5", X"002C", X"FA67", X"FAE7", X"FAC7", X"FD9B", X"FF1A", X"FEA1", X"FFE3", X"0298", X"0268", X"00E0", X"0173", X"00F4", X"01A2", X"FFE5", X"00B4", X"FF95", X"FCBC", X"FE56", X"FD13", X"FEC8", X"FDD4", X"FE4B", X"FEF0", X"00E2", X"0348", X"0045", X"0191", X"FFAC", X"FC3C", X"FD78", X"FC59", X"FD4E", X"FC58", X"FE2D", X"00E4", X"0295", X"0322", X"0250", X"036E", X"01DF", X"02C1", X"0154", X"02E1", X"0174", X"FE29", X"FE87", X"FEBE", X"FE61", X"FD62", X"FE14", X"FE22", X"011E", X"01E8", X"0123", X"FFA1", X"0030", X"FD5E", X"FC31", X"FAFA", X"FC0D", X"FC8E", X"FB00", X"FE4B", X"FF34", X"FEC5", X"002A", X"FD19", X"FD2E", X"FEDC", X"0146", X"01F8", X"02A7", X"036E", X"0433", X"042D", X"019A", X"003E", X"021B", X"FAEB", X"FD31", X"FD88", X"003E", X"00E3", X"0024", X"014B", X"009C", X"FC08", X"FC59", X"FB17", X"FB3A", X"F86C", X"F90D", X"FB3B", X"F8E1", X"F94B", X"FA81", X"FDAA", X"FF83", X"00F3", X"033A", X"062A", X"07CA", X"0824", X"08DD", X"0589", X"050A", X"0117", X"FDCC", X"FDA7", X"FEFC", X"009B", X"FF5E", X"FF3C", X"021F", X"0013", X"0125", X"002F", X"FFF1", X"FFD8", X"FF19", X"FF24", X"007A", X"FFA6", X"0095", X"0143", X"FE18", X"0089", X"00A6", X"03F8", X"03C2", X"044E", X"0438", X"037C", X"014E", X"0062", X"FEB1", X"0063", X"FEA9", X"0070", X"000F", X"012F", X"0152", X"005F", X"001F", X"004F", X"0203", X"FF73", X"FF07", X"FF36", X"FF70", X"FDB7", X"FCA2", X"0114", X"FD9B", X"FF7C", X"FB93", X"FD3B", X"FF96", X"FFCB", X"FFEF", X"014F", X"FFF3", X"FFE8", X"FE5F", X"FFDF", X"008F"),
        (X"FE4D", X"0071", X"FF79", X"0015", X"FFE3", X"FECB", X"007D", X"004D", X"FFF8", X"0003", X"0104", X"FFFB", X"FF2A", X"FEAD", X"0026", X"FFCC", X"FFC4", X"FF44", X"FF25", X"FFF0", X"010E", X"0167", X"FFF7", X"0065", X"FFD1", X"011D", X"0087", X"0012", X"0119", X"019F", X"0145", X"003A", X"FFDF", X"FE74", X"FCA1", X"FBF5", X"FBB8", X"FB81", X"FBB6", X"F935", X"FA48", X"FA09", X"FF22", X"FAF7", X"FB44", X"FAEE", X"FA72", X"FB96", X"FB8F", X"FCDC", X"FBE8", X"FCFD", X"FE29", X"00C7", X"008B", X"0149", X"FED1", X"FFC8", X"FFFB", X"FD98", X"FC83", X"FCF3", X"FCAD", X"F939", X"F7AD", X"F671", X"F5CB", X"F512", X"F282", X"F901", X"FA7D", X"F71D", X"FC40", X"FBF9", X"F8EA", X"F7AC", X"F767", X"FA0B", X"FA77", X"FC43", X"FBE9", X"FE27", X"006A", X"013D", X"0044", X"0066", X"00A7", X"FD8F", X"FCB9", X"FB33", X"FA10", X"F5DA", X"F6F1", X"F6BC", X"F7B4", X"F672", X"F4D4", X"F3E4", X"F573", X"F871", X"F81E", X"FA3C", X"FA95", X"FB43", X"F7F2", X"FB81", X"FCE2", X"FCA8", X"FBDF", X"FBCE", X"FDCE", X"011A", X"FF74", X"FF9A", X"0078", X"FF25", X"FFE6", X"00FF", X"FEC8", X"FCC2", X"FA62", X"FAE0", X"F755", X"F6E9", X"F7DF", X"F96A", X"F7B4", X"F78C", X"F7BB", X"F839", X"F8E3", X"FF5E", X"0122", X"013F", X"02A0", X"01FB", X"0079", X"FB03", X"FB88", X"FDFA", X"0089", X"000D", X"FEA5", X"FECA", X"FFD1", X"0299", X"025B", X"FEBE", X"019D", X"00B8", X"FD76", X"FDB3", X"FCEF", X"FE1F", X"FE68", X"FFEF", X"FEAA", X"FD25", X"FE61", X"FCFB", X"FE03", X"FF21", X"FFF1", X"0325", X"018B", X"FCD3", X"FB89", X"FF55", X"001D", X"FEC9", X"0171", X"02FA", X"00B8", X"028B", X"0245", X"002E", X"FFF8", X"0084", X"FF45", X"FF86", X"0054", X"0034", X"FF7A", X"0081", X"FEBC", X"007F", X"FF8E", X"FEE8", X"FDD4", X"FFEB", X"FE94", X"FD79", X"FF7D", X"FAF5", X"FF1A", X"FE34", X"009C", X"FC76", X"03D8", X"06AF", X"02D9", X"0264", X"FFD0", X"005D", X"FFBA", X"FF91", X"01BB", X"FFFD", X"FDFE", X"FF69", X"FE5E", X"FD22", X"FDD7", X"FFFE", X"00C7", X"0027", X"0067", X"FF88", X"FEE9", X"FEF2", X"FD1B", X"FCCE", X"0110", X"FE3B", X"00CF", X"FFA1", X"02C3", X"02CC", X"0195", X"0035", X"FF00", X"0080", X"FFCD", X"FF48", X"FF05", X"00BD", X"FF26", X"FDAE", X"FDEA", X"FF21", X"FC92", X"00E5", X"0285", X"FE3E", X"FF00", X"FF27", X"FED9", X"FEA0", X"FC83", X"FE9F", X"FBF5", X"FD41", X"00B7", X"0448", X"020A", X"0331", X"FD06", X"FD38", X"FE28", X"FF99", X"FF80", X"00A4", X"0072", X"003E", X"00AE", X"FE66", X"FE5C", X"FF3C", X"01DA", X"01C3", X"0333", X"002F", X"FEE3", X"FEDC", X"FFAE", X"FAFC", X"FA49", X"F935", X"F90F", X"0019", X"022F", X"0560", X"01BA", X"02A5", X"FC9C", X"FDEC", X"FE52", X"FF64", X"FFA1", X"0077", X"FFF2", X"FFD2", X"0102", X"FBF8", X"FBD1", X"02B3", X"0640", X"0346", X"0382", X"0321", X"00CC", X"00EF", X"FF5A", X"F7F1", X"F6C8", X"F80B", X"F757", X"FD44", X"0146", X"02C7", X"0149", X"007A", X"FDBE", X"FDA0", X"0048", X"01A1", X"0217", X"018F", X"02D9", X"02D3", X"005F", X"FA96", X"FE95", X"077C", X"0813", X"06B7", X"04D1", X"02F8", X"0377", X"024A", X"FF73", X"F79B", X"F25A", X"F655", X"F94E", X"FEDF", X"0213", X"0256", X"03CF", X"FF74", X"FE81", X"FFA8", X"0034", X"010D", X"021B", X"00CA", X"02E8", X"01D4", X"FEA2", X"FA69", X"0112", X"08A2", X"0802", X"076E", X"0545", X"023B", X"0288", X"0299", X"01B0", X"FB95", X"F441", X"FAAD", X"FF9F", X"FFD8", X"FFB7", X"01BB", X"02EA", X"FF85", X"037D", X"013C", X"0249", X"024F", X"0144", X"00D0", X"01D2", X"01F7", X"FBED", X"FC43", X"042F", X"062B", X"03E1", X"0535", X"04A4", X"03EB", X"04BC", X"04CA", X"020D", X"F9C9", X"FAEB", X"FACE", X"FB24", X"FCD5", X"FDFC", X"0180", X"01AB", X"0176", X"05BE", X"032C", X"02C5", X"02EA", X"02B1", X"0287", X"001B", X"FF31", X"FC9B", X"FE87", X"02CF", X"02C9", X"04F2", X"0638", X"0629", X"08A3", X"0624", X"0390", X"01B4", X"FD27", X"FC72", X"FBAD", X"FA93", X"FD40", X"FF39", X"FFDE", X"0241", X"0240", X"0735", X"04FE", X"039C", X"026E", X"015B", X"FFFD", X"FF08", X"FF53", X"FE15", X"FD31", X"FFF6", X"03B6", X"047B", X"0459", X"0693", X"0687", X"0422", X"039C", X"01B8", X"FEDE", X"F84C", X"FA14", X"FF3B", X"FF0C", X"02A5", X"FF39", X"FDF7", X"FE52", X"061A", X"052A", X"048B", X"064A", X"04EC", X"0066", X"FD1C", X"FD4A", X"FCD6", X"FF15", X"010B", X"02F1", X"0313", X"0768", X"075F", X"041A", X"0311", X"0073", X"013E", X"FD54", X"F936", X"F74F", X"FB61", X"FFDE", X"FFC2", X"FF29", X"FEB6", X"FD66", X"01FE", X"00A2", X"0080", X"0373", X"0320", X"0202", X"0144", X"FF60", X"008C", X"031E", X"03D6", X"05DC", X"0415", X"0556", X"030D", X"00DE", X"0132", X"0178", X"FEA9", X"FC7C", X"FA43", X"FC2C", X"FD5C", X"FEC8", X"01F3", X"FF43", X"0025", X"FE3B", X"007D", X"FEAD", X"FE18", X"FF98", X"023C", X"0317", X"00EF", X"0212", X"0193", X"032D", X"045C", X"04C2", X"00DD", X"FED4", X"FF6E", X"FD55", X"0015", X"FF08", X"FA89", X"F992", X"F858", X"FA9D", X"FF54", X"0163", X"00FC", X"FE59", X"0156", X"0081", X"004A", X"FDC9", X"FBEB", X"FD77", X"FE64", X"FC1C", X"FB95", X"FC55", X"F9A2", X"FCDE", X"FF59", X"FD26", X"FC8F", X"FAFD", X"FAE2", X"FBB4", X"FB42", X"FB86", X"F57E", X"F5AC", X"F87C", X"FB11", X"FDFD", X"0243", X"0112", X"FDD1", X"FFA8", X"FD7F", X"FB34", X"F94F", X"FA2D", X"F850", X"F87B", X"F92A", X"F89F", X"F8D0", X"F815", X"F946", X"F976", X"FA12", X"FB83", X"FAE2", X"F7DA", X"F8A3", X"F99F", X"F8EE", X"F59A", X"F656", X"FBB5", X"FB54", X"FD2C", X"0079", X"016D", X"FFF8", X"FB47", X"F9F0", X"FB62", X"FD01", X"FA34", X"FB19", X"FAAF", X"FB4A", X"FB32", X"F9A4", X"F8D5", X"F73D", X"F95E", X"FA4D", X"FBD4", X"F809", X"F89C", X"FA4B", X"FA0B", X"F84F", X"F6AF", X"F842", X"FDEB", X"FDEF", X"FE97", X"FF70", X"00A6", X"0149", X"FC35", X"F947", X"FD3B", X"0104", X"FF54", X"FE17", X"FF5F", X"FDBF", X"FFDB", X"FC02", X"FB34", X"FABA", X"FACB", X"FC04", X"FAC2", X"FB6C", X"FB5A", X"FCFC", X"FBCC", X"FBCC", X"FAC4", X"FB2E", X"FF2B", X"FDD9", X"FE58", X"FED8", X"FFC4", X"012B", X"FC15", X"FAD6", X"0046", X"01AE", X"03D7", X"0208", X"002F", X"FF1A", X"00DD", X"FE05", X"FCF0", X"FD26", X"FD3F", X"FAD1", X"FC01", X"FD37", X"FCE9", X"FE37", X"FD17", X"FED9", X"FF08", X"FC8F", X"FE8D", X"FED7", X"FF06", X"00BF", X"FF66", X"FFF6", X"FEB7", X"FF1A", X"047D", X"084E", X"042E", X"03F3", X"01D1", X"FF20", X"FE75", X"FE75", X"FB00", X"FB12", X"FA11", X"FAE0", X"FA7A", X"FC4B", X"FBD2", X"FDD9", X"FF6C", X"0339", X"0121", X"FEB4", X"FB61", X"FC01", X"FDB6", X"0059", X"0104", X"0078", X"FF85", X"025E", X"054B", X"06EB", X"01D8", X"022F", X"0050", X"FF7F", X"FDD2", X"FFAB", X"FE8F", X"FC08", X"FC57", X"FEA7", X"FB77", X"FBC8", X"FE4E", X"FF2E", X"0382", X"0441", X"FF06", X"0142", X"FD60", X"FE42", X"FE46", X"0091", X"0003", X"FF2A", X"FFA9", X"FF9D", X"0141", X"022A", X"048A", X"062F", X"0584", X"0570", X"03C8", X"00E3", X"FF69", X"01B8", X"0425", X"0295", X"0240", X"0391", X"0363", X"028D", X"01F4", X"01B9", X"003F", X"0089", X"0046", X"011C", X"0137", X"FE42", X"FF20", X"FF11", X"00E2", X"0168", X"FF8E", X"FFB6", X"FFE3", X"0092", X"0205", X"0275", X"0070", X"FF6A", X"0163", X"02EB", X"067D", X"05E8", X"05F6", X"05AA", X"03C9", X"03DB", X"0391", X"0401", X"042C", X"014F", X"FFE2", X"FE70", X"0036", X"0018"),
        (X"017F", X"FF3C", X"002B", X"0247", X"0028", X"000A", X"FF43", X"FFC6", X"0052", X"FF9D", X"FF7B", X"FF0A", X"FD12", X"0022", X"00BC", X"FF6B", X"FF23", X"0061", X"FED0", X"FF9A", X"FF23", X"007E", X"FF21", X"000F", X"000A", X"FE25", X"0042", X"FFA7", X"FFBD", X"0232", X"0028", X"FF37", X"FF76", X"0083", X"FEA9", X"FEC3", X"FCD7", X"FB3E", X"F9F5", X"FA01", X"F90E", X"FA5E", X"FCCE", X"FD8D", X"FD35", X"FB9C", X"FB70", X"FCE9", X"FA3E", X"FE08", X"FCDB", X"FE31", X"FF78", X"00B4", X"FF5C", X"FF86", X"FF84", X"0014", X"FECF", X"FE13", X"FCF4", X"FF75", X"FBBD", X"F8B0", X"F980", X"FB35", X"FA28", X"FCAF", X"FD08", X"FBCC", X"FAF3", X"FCD9", X"FC6B", X"FB68", X"FA96", X"F962", X"FC28", X"FC3B", X"FC4A", X"FBA7", X"FF9F", X"FECA", X"FFC3", X"FE6F", X"FECA", X"0011", X"FF6D", X"FC6F", X"FC98", X"FEF6", X"FE9D", X"0012", X"FE45", X"FEC6", X"FF8C", X"000E", X"FF7A", X"FE66", X"FB48", X"FB45", X"FBA8", X"FCD6", X"FDB9", X"FEE1", X"FE5A", X"FD2A", X"FC72", X"FDF3", X"FE98", X"FFEF", X"0065", X"FFE5", X"FF55", X"FFF2", X"FE2C", X"016E", X"FDC2", X"FFC2", X"00F6", X"0272", X"0134", X"FF54", X"FECA", X"017A", X"00E9", X"010B", X"027B", X"000E", X"FF37", X"FF4D", X"0091", X"FF77", X"FE7F", X"FFA8", X"FCE9", X"FBD1", X"FF7B", X"00CD", X"0274", X"FFF8", X"006B", X"0079", X"0027", X"02C4", X"0204", X"00EC", X"0039", X"FF3D", X"FEDB", X"FF79", X"FD2D", X"FDA6", X"FF89", X"FDA3", X"FCB1", X"FF45", X"025D", X"0262", X"006F", X"01D0", X"006C", X"0109", X"FF3C", X"FDF1", X"FEEF", X"0319", X"FEFA", X"0221", X"0088", X"0097", X"FDD1", X"041B", X"019B", X"023D", X"0008", X"FF09", X"FF37", X"FE39", X"FE6A", X"FC39", X"FBDD", X"FBA6", X"FD47", X"001E", X"0108", X"01DE", X"002F", X"FF8D", X"FE9E", X"0039", X"FFAD", X"FF73", X"0238", X"0080", X"00B4", X"038B", X"00B0", X"0042", X"0184", X"076D", X"07B8", X"03A0", X"FFAF", X"FEA3", X"006D", X"FFAE", X"FE26", X"FF6F", X"FBF0", X"FBF1", X"FC6E", X"FE6A", X"FFF9", X"0008", X"01C7", X"0186", X"0018", X"FFCF", X"02CD", X"03A2", X"01FB", X"0126", X"021D", X"01B7", X"FFDD", X"02CC", X"02CB", X"079F", X"0745", X"03A8", X"014C", X"0149", X"00D4", X"0063", X"010F", X"FCF4", X"FD2A", X"FDE1", X"FCE5", X"00EF", X"034B", X"0555", X"043C", X"04C4", X"0138", X"027C", X"063C", X"04FA", X"0872", X"062D", X"0421", X"02C2", X"0129", X"039F", X"069E", X"0732", X"051E", X"047C", X"00D7", X"02D3", X"01B8", X"0129", X"005A", X"FC04", X"F9F9", X"FC41", X"00C6", X"06C0", X"07CB", X"06B6", X"04E4", X"05CF", X"0320", X"03E4", X"0856", X"06FA", X"0846", X"07BA", X"0528", X"FF76", X"0363", X"04B6", X"07F2", X"06D0", X"034B", X"0167", X"0259", X"0085", X"FE7D", X"FD72", X"FC08", X"F9E5", X"FA98", X"0069", X"088B", X"0AF6", X"04B3", X"0212", X"04B3", X"04F8", X"0152", X"00A8", X"04AC", X"03C8", X"057D", X"0463", X"0509", X"0007", X"00D6", X"03F3", X"0504", X"02A1", X"0225", X"0174", X"FD7A", X"FD70", X"FCE7", X"FBEA", X"F94B", X"FAD8", X"FD54", X"04EB", X"0B71", X"05EA", X"FE0B", X"FC86", X"005E", X"011B", X"FF19", X"FF0D", X"FEFD", X"FFB1", X"02A9", X"0741", X"0414", X"00D2", X"0038", X"0056", X"012C", X"FEEA", X"FD32", X"FBF1", X"FAD8", X"FA11", X"FAA3", X"FB4E", X"FA43", X"FDFB", X"0282", X"07FC", X"0926", X"0163", X"FEBE", X"FC35", X"FF6B", X"00B8", X"FF05", X"FEAF", X"FAFB", X"F8E1", X"FEDB", X"0621", X"072E", X"02A6", X"0032", X"FEA7", X"FE9C", X"FE31", X"F6D2", X"F7CA", X"F789", X"F982", X"FAFD", X"FF25", X"FDEC", X"006C", X"05C6", X"0800", X"06DA", X"034E", X"FF6E", X"FEB1", X"0190", X"FF58", X"000C", X"FCFF", X"F9E8", X"F8E1", X"FCC0", X"0655", X"07A6", X"02F9", X"FE2E", X"FBC9", X"0124", X"FDA9", X"F5BD", X"F777", X"F869", X"FA1A", X"FD82", X"000F", X"015C", X"02D5", X"06C1", X"095C", X"065C", X"024C", X"FFEA", X"FF80", X"FFDD", X"FEBE", X"FE4E", X"FD8B", X"FC79", X"FA7E", X"FBBD", X"031A", X"08F9", X"02DA", X"00C9", X"FE3E", X"FECB", X"012D", X"F9D5", X"FB43", X"FBB7", X"FC2B", X"FE85", X"0198", X"00CC", X"012F", X"0508", X"083A", X"094F", X"0533", X"FF5F", X"FEAA", X"FD8B", X"FFB3", X"FDDE", X"FE4A", X"FCB9", X"FDCE", X"00DC", X"0385", X"06B4", X"0236", X"0032", X"014D", X"0360", X"053F", X"00D1", X"FC26", X"FCC0", X"FDD1", X"FD22", X"0174", X"FF51", X"FF9C", X"0510", X"0976", X"09D4", X"0465", X"000C", X"FEAD", X"FDF6", X"FE7A", X"FE96", X"004B", X"FE37", X"0263", X"0323", X"0474", X"089C", X"02D0", X"0019", X"FFA5", X"033B", X"044D", X"03CC", X"FE0C", X"FFBA", X"FF2F", X"FF8C", X"FF1B", X"FFAB", X"FFA6", X"0465", X"0AC3", X"084B", X"0114", X"FE96", X"FCC0", X"FD44", X"FEDB", X"FED7", X"0035", X"0166", X"01A0", X"04BF", X"037E", X"0599", X"0071", X"FF99", X"00C8", X"00E4", X"0109", X"024B", X"0400", X"04C0", X"00AA", X"00BF", X"FD99", X"FCD2", X"FFD2", X"04E1", X"0B70", X"0462", X"FD3B", X"FB8D", X"FCE5", X"FD5A", X"FE67", X"FEB0", X"FE80", X"0363", X"0486", X"036C", X"0116", X"028C", X"01DE", X"00CF", X"022D", X"FD35", X"FF2B", X"FF2F", X"02BA", X"02E6", X"0270", X"FFBB", X"0172", X"00C4", X"00E7", X"0746", X"09BA", X"FFD0", X"FAC2", X"F9DD", X"FD48", X"FF24", X"FE9A", X"FF89", X"013C", X"02B8", X"03A0", X"FE05", X"0190", X"03DA", X"0238", X"FFCD", X"FFCF", X"FDD1", X"00F9", X"FF0C", X"00AF", X"04CF", X"0335", X"0361", X"030A", X"04E4", X"05D7", X"0785", X"036F", X"FDF8", X"F8A6", X"FA24", X"FD0D", X"FE41", X"FF71", X"FF8E", X"0214", X"034E", X"014B", X"0061", X"FED2", X"00E2", X"FE25", X"FFC4", X"031C", X"026F", X"04F7", X"FDD3", X"0006", X"00D8", X"0316", X"012C", X"029A", X"0500", X"038B", X"0266", X"FF63", X"FBCB", X"FA7C", X"FA56", X"FC97", X"FE3A", X"FDC4", X"FFA9", X"FF9C", X"0057", X"00BD", X"FD90", X"FD5F", X"FE35", X"FF03", X"FFDE", X"FF5E", X"0536", X"0419", X"0196", X"FF3B", X"01E9", X"024F", X"0407", X"0373", X"0400", X"02E3", X"0028", X"FAA1", X"FB96", X"FB21", X"FAF1", X"FD3C", X"FDEA", X"FFF6", X"FF42", X"FF07", X"00E6", X"009E", X"FF34", X"FD4D", X"FC2F", X"FFF7", X"FFA7", X"00D3", X"028F", X"0147", X"04A5", X"018C", X"0203", X"0312", X"0360", X"03E3", X"0264", X"004D", X"FD25", X"FCE2", X"FBC3", X"FDF5", X"FDC3", X"FDFE", X"FFC5", X"01B9", X"0067", X"FE75", X"FE4A", X"FCEF", X"FC15", X"FE89", X"0024", X"001C", X"FFBE", X"0035", X"FF74", X"FE3C", X"00A8", X"0181", X"0133", X"031D", X"0424", X"01C6", X"FF34", X"FDBB", X"FC53", X"FD70", X"00B7", X"FE98", X"FE61", X"FBC3", X"FDB4", X"FE4B", X"FE0A", X"FD91", X"FB02", X"FD2D", X"0229", X"0409", X"021B", X"00F4", X"00C4", X"0033", X"004A", X"FCDE", X"00A2", X"FF7A", X"021A", X"04D2", X"0568", X"04C0", X"0226", X"FE1E", X"FCE3", X"FB8F", X"FE99", X"FFC7", X"FF11", X"FD50", X"FC79", X"FBBD", X"F9B6", X"F8E8", X"F6E8", X"FB7E", X"FD63", X"0128", X"0271", X"010E", X"0068", X"FFD9", X"FE76", X"0059", X"FF9E", X"FC2F", X"FF64", X"0244", X"0037", X"FF1E", X"FF8B", X"FB84", X"FA4F", X"FA0B", X"F6A8", X"F8E2", X"F8C7", X"F7FC", X"F730", X"F6AD", X"F6D1", X"F71C", X"FB0C", X"FDA9", X"FDA5", X"0070", X"00A8", X"FFC7", X"0005", X"017F", X"009C", X"002E", X"FF48", X"0269", X"011A", X"010C", X"039C", X"048D", X"01DC", X"0285", X"0224", X"069F", X"0093", X"030F", X"0755", X"0807", X"0186", X"004E", X"FCFA", X"FE04", X"FF9A", X"0255", X"FFEB", X"FE14", X"FF4C", X"0089"),
        (X"0088", X"FFD9", X"008A", X"FF51", X"027D", X"FFA9", X"FF9B", X"0090", X"017F", X"FFC4", X"FF54", X"FFD9", X"FF03", X"FF6B", X"FFF9", X"00CD", X"00C9", X"00BC", X"0048", X"FEC2", X"0140", X"0063", X"FF80", X"FF50", X"FF36", X"00DD", X"0026", X"0186", X"0014", X"FF6A", X"0077", X"FF71", X"0072", X"FF26", X"0042", X"FF67", X"014F", X"FF45", X"0263", X"FE5D", X"FF6A", X"FF8C", X"FEBC", X"FDAB", X"0125", X"00F2", X"0158", X"01BE", X"0164", X"01E4", X"005B", X"005A", X"FF8B", X"00B0", X"FFB1", X"00F0", X"0053", X"FFDD", X"FE88", X"FC90", X"FE12", X"0088", X"029D", X"02BC", X"030A", X"05F1", X"0507", X"078A", X"0403", X"050D", X"02DD", X"FE98", X"FE36", X"FF54", X"0008", X"0107", X"024C", X"02AF", X"00B1", X"0138", X"02AE", X"0073", X"FFE5", X"0065", X"FFC3", X"FF11", X"FE4D", X"FB51", X"FF88", X"FE5F", X"FEC6", X"0086", X"FFC0", X"039A", X"0299", X"02E2", X"01F0", X"017A", X"00CB", X"FD85", X"FD34", X"FE02", X"FDE6", X"FF28", X"0064", X"034E", X"060E", X"076D", X"0684", X"0261", X"02A4", X"FF65", X"0051", X"0105", X"FC30", X"FBE2", X"003F", X"FDBB", X"FE88", X"FE39", X"FF56", X"FF6E", X"0092", X"0066", X"001F", X"FFE0", X"FFE8", X"FE1F", X"FE61", X"00E3", X"FE8D", X"FF99", X"0270", X"00D6", X"0210", X"03DD", X"0400", X"0419", X"01B8", X"02CB", X"FF1B", X"FFB1", X"FDEA", X"FB9E", X"FF8E", X"FE29", X"FE1C", X"00A2", X"0255", X"01AD", X"044C", X"0487", X"062C", X"01E1", X"0226", X"01F0", X"01B1", X"0388", X"00B7", X"0180", X"01A1", X"01B5", X"0073", X"0136", X"0288", X"076D", X"00AE", X"0153", X"0157", X"FDDD", X"FE3D", X"FD05", X"FFA0", X"00A2", X"00C9", X"01A6", X"0423", X"031C", X"010C", X"02A0", X"0534", X"0650", X"0419", X"051A", X"0249", X"0132", X"FFD8", X"01BD", X"00B5", X"002C", X"FE95", X"FF29", X"0169", X"03EE", X"00FE", X"021A", X"FEC9", X"FD5C", X"FF72", X"FA49", X"014A", X"0038", X"013B", X"0050", X"00AA", X"FF6D", X"018F", X"016D", X"02E5", X"03C7", X"009D", X"017E", X"014E", X"FE17", X"FDBB", X"FBBD", X"FD36", X"0045", X"FFB9", X"FE22", X"FF7E", X"FFA7", X"0133", X"FF7C", X"FDFE", X"FE2B", X"FF4A", X"FBBC", X"0032", X"FFAD", X"00DE", X"0026", X"FEA0", X"FFC2", X"0134", X"0160", X"0125", X"005D", X"FC01", X"FB1A", X"F954", X"FB95", X"F9BA", X"FB5B", X"FA94", X"FD83", X"FED6", X"FEF4", X"FAE0", X"FD1D", X"FE3C", X"FF80", X"FE53", X"FB51", X"FDA7", X"FBE4", X"FEC3", X"FF5E", X"FF7C", X"FC89", X"FF9E", X"FFFB", X"029A", X"02E5", X"0161", X"FD00", X"FA51", X"F8CA", X"F96E", X"FA0A", X"FBB6", X"FB5F", X"FB15", X"FC8F", X"FB5C", X"FCA9", X"F5F9", X"F7BF", X"FA63", X"FBB7", X"FDF2", X"FCEC", X"FAC5", X"FB25", X"FDC7", X"0066", X"01C4", X"002D", X"FF9B", X"0068", X"029E", X"0460", X"037F", X"FBE5", X"FA86", X"F714", X"FB2E", X"FB40", X"FAEC", X"FD17", X"FACA", X"FABD", X"FD47", X"FBFA", X"F62A", X"F4CD", X"F849", X"FDB2", X"FF1A", X"FAB8", X"F865", X"F969", X"FCAC", X"01E8", X"011A", X"FFBA", X"0009", X"FD62", X"0100", X"06C6", X"FFE6", X"F9F3", X"F72A", X"F6B5", X"FA6D", X"FD13", X"FD90", X"FDEE", X"FE7F", X"FE3D", X"01A9", X"FE58", X"F9D0", X"F703", X"F9B5", X"FBB1", X"FFCB", X"FBDE", X"FAC8", X"FCF4", X"FF28", X"001E", X"FE76", X"FC72", X"FCEA", X"FE08", X"03B2", X"0532", X"0101", X"FD64", X"FA7F", X"FCF9", X"FF90", X"FFF6", X"FC84", X"FFD4", X"0165", X"01F7", X"038A", X"03E1", X"02A6", X"FF6A", X"FDD7", X"FDB3", X"FFBA", X"FE0B", X"FACE", X"FF02", X"00B3", X"FF88", X"FD2A", X"FAFD", X"FC3B", X"FCDB", X"03A8", X"07AE", X"0707", X"00E0", X"0063", X"0144", X"0410", X"03F9", X"0187", X"01A2", X"0127", X"02D3", X"01E4", X"0261", X"0145", X"FFD7", X"042F", X"0366", X"FEC4", X"FE7F", X"FACA", X"FEED", X"00CF", X"FC96", X"FEF1", X"FDC3", X"FD85", X"0070", X"04DA", X"09A9", X"0771", X"02B0", X"00E3", X"02C8", X"0604", X"0424", X"002C", X"FFBB", X"FF3C", X"FF25", X"FC5D", X"FD55", X"FB0C", X"030D", X"03F7", X"013E", X"FFA7", X"FF46", X"FDAB", X"0157", X"014E", X"000C", X"FDCD", X"FD31", X"FDE4", X"0202", X"0876", X"0632", X"07E0", X"045C", X"024A", X"0434", X"05D5", X"05C2", X"017C", X"00AB", X"FF09", X"FD79", X"FD02", X"FAA7", X"FB7A", X"0577", X"04CF", X"02BF", X"FEB3", X"FF6D", X"FD86", X"01DC", X"FEF5", X"FE72", X"FE9C", X"FEE9", X"0010", X"040B", X"07D2", X"0860", X"0788", X"04B1", X"0191", X"03BE", X"04F9", X"03F2", X"01C2", X"FF58", X"00C7", X"FF9D", X"0023", X"FE53", X"FF18", X"0A0C", X"0556", X"015A", X"FFCA", X"FE50", X"FF47", X"FFEC", X"FE0A", X"FE15", X"00EB", X"FF41", X"01AB", X"0566", X"0801", X"094A", X"0820", X"025B", X"00F0", X"045A", X"02B8", X"0214", X"0448", X"0405", X"01F3", X"0014", X"FE36", X"FE6C", X"0038", X"03A4", X"0127", X"FE73", X"FE68", X"FF61", X"FDC8", X"FDE1", X"FEDB", X"FDAF", X"FF6B", X"FE0D", X"FCBF", X"00A1", X"0246", X"02D3", X"02C9", X"FF77", X"FEF2", X"0302", X"02B7", X"025B", X"03D0", X"02DC", X"FF54", X"FD67", X"FE61", X"0192", X"02EA", X"0325", X"FE51", X"0036", X"FF7B", X"FA47", X"FEC8", X"FEEC", X"0005", X"FF9F", X"FE28", X"FB74", X"FBF0", X"FD17", X"FFAB", X"0021", X"00F6", X"FE6B", X"009F", X"01DE", X"0405", X"03A2", X"032A", X"FFAD", X"FE75", X"FFBA", X"FE52", X"0232", X"00E6", X"FEAE", X"FE9B", X"FE14", X"022C", X"FD3C", X"FDAA", X"FD1B", X"0069", X"FE9E", X"FD18", X"FE69", X"FAB7", X"FA93", X"FDBA", X"FD53", X"FE75", X"0086", X"015B", X"02C6", X"02EA", X"FFEA", X"016E", X"01C9", X"0267", X"00CC", X"009C", X"04A8", X"0184", X"0158", X"FE6B", X"FEE1", X"FF7F", X"002D", X"FF8A", X"FE64", X"FE6C", X"FEA4", X"FC5A", X"FF57", X"FC55", X"FCF5", X"FBB3", X"FE32", X"0090", X"01A9", X"0222", X"006F", X"00B7", X"039E", X"02C1", X"0198", X"00EE", X"FD38", X"02D7", X"06F5", X"0403", X"00BA", X"FD03", X"00B2", X"FE5C", X"FF57", X"01D8", X"0067", X"FFBC", X"FD08", X"FE4D", X"FE45", X"FF18", X"FF0A", X"00D9", X"00D3", X"0204", X"0286", X"0149", X"FE83", X"012D", X"FFBC", X"0093", X"0090", X"035F", X"00F8", X"04DA", X"07ED", X"05FA", X"017E", X"FC69", X"000D", X"009F", X"FF92", X"FBFE", X"006B", X"FE1C", X"FA7D", X"FBAC", X"FBD8", X"001E", X"FF38", X"0012", X"011A", X"00B3", X"036C", X"FFA6", X"FF74", X"00A2", X"0043", X"0168", X"0387", X"05FF", X"0764", X"0829", X"08BB", X"0423", X"FFF0", X"FBDA", X"005C", X"FF2B", X"FFC7", X"FC45", X"F8E7", X"F791", X"F76C", X"F7F2", X"FB77", X"FF1E", X"0150", X"00C6", X"00A8", X"01B4", X"FFED", X"FF5E", X"0164", X"02E6", X"01CC", X"0374", X"058B", X"078A", X"05F6", X"06C3", X"0631", X"0210", X"00FE", X"FDFE", X"015A", X"016C", X"FEFE", X"FFD8", X"FC75", X"FAE1", X"FD1A", X"FE32", X"FB72", X"FAC9", X"FBC7", X"FEB1", X"FD96", X"FAD5", X"FCBD", X"FFDE", X"0168", X"000E", X"FE93", X"002C", X"FD85", X"016D", X"0317", X"002A", X"02EA", X"FE62", X"002C", X"FFB9", X"FE64", X"FFBD", X"0049", X"FEBD", X"020F", X"0502", X"03CC", X"0463", X"0481", X"03F8", X"03AB", X"02C8", X"FF16", X"FFD0", X"FD73", X"FFB7", X"FD94", X"FB91", X"FDF5", X"FDAC", X"FBA1", X"00A4", X"0344", X"FE65", X"02C8", X"0059", X"FFAE", X"0074", X"0030", X"01B4", X"FFD1", X"FF8A", X"FF81", X"FFEF", X"FE13", X"026E", X"FFBB", X"FE82", X"FEAD", X"FD0F", X"000D", X"0009", X"FC18", X"00A3", X"0143", X"FDDB", X"FBFA", X"FDF7", X"FCC6", X"FFBE", X"FE38", X"0109", X"FDD1", X"0018", X"FF48", X"0007", X"FFD3"),
        (X"00C0", X"FED1", X"01B7", X"FF6D", X"00D6", X"00A5", X"FF3B", X"00B0", X"FE86", X"FFEF", X"0054", X"FFB0", X"FE23", X"FDE0", X"0078", X"FFB1", X"003B", X"0030", X"FF6C", X"00CE", X"FEB9", X"FF5A", X"00A4", X"005F", X"FF57", X"003F", X"FFD5", X"0087", X"0124", X"0055", X"FF55", X"0024", X"0165", X"0088", X"FD4C", X"FBF3", X"FB42", X"FCDB", X"FB73", X"FB46", X"F9E2", X"FC10", X"0057", X"01EC", X"0233", X"FE2D", X"FAE6", X"FB57", X"FBFB", X"FCB6", X"FEE7", X"FE30", X"0114", X"00AB", X"FF1A", X"0095", X"FF90", X"0080", X"FFE0", X"FD35", X"FDF6", X"FEA4", X"FB23", X"F849", X"FAD8", X"00BA", X"FE91", X"FF6D", X"FEA5", X"007D", X"00B6", X"035F", X"0402", X"0318", X"01A9", X"FE6B", X"FC5B", X"FCB8", X"FADF", X"FD31", X"011F", X"0264", X"010C", X"0102", X"FEF1", X"FED3", X"00B2", X"FF2C", X"FED3", X"0169", X"FC4C", X"FE7D", X"FF35", X"0024", X"00D4", X"FFBC", X"0481", X"04D8", X"0403", X"04AB", X"03FB", X"01ED", X"FE3C", X"FF1D", X"FDCC", X"FE1B", X"F88B", X"F6BD", X"FADF", X"FFA2", X"FDAE", X"FF79", X"FF9C", X"0173", X"01A4", X"036F", X"021D", X"02EF", X"00A7", X"00BC", X"01AB", X"01E7", X"02F6", X"0069", X"0285", X"0396", X"03AA", X"028D", X"00F7", X"00DE", X"010A", X"002D", X"FD5F", X"FA9B", X"F826", X"F6A4", X"F5CC", X"F9FC", X"FB33", X"FD99", X"FFCB", X"FF88", X"01F2", X"025F", X"07DC", X"0662", X"0158", X"01A8", X"0148", X"FF5E", X"0060", X"0043", X"0163", X"0196", X"030A", X"0430", X"032D", X"01FB", X"005B", X"FFDC", X"FDB9", X"FE41", X"FC5B", X"F980", X"F8EF", X"F78C", X"FD5B", X"FD93", X"002A", X"FF17", X"FF1E", X"071F", X"07A6", X"0532", X"044A", X"0017", X"0020", X"FFCD", X"008B", X"FFC3", X"01B8", X"013C", X"01A5", X"010B", X"0314", X"00B8", X"017B", X"FF64", X"FE9A", X"FED1", X"FD72", X"FAA4", X"F90E", X"F680", X"FC8E", X"FE71", X"005E", X"0149", X"033E", X"0801", X"09B1", X"05A7", X"024F", X"FE72", X"FE28", X"FC5A", X"FF56", X"FFE7", X"0265", X"029D", X"0266", X"FFED", X"FE57", X"FEE8", X"002D", X"010E", X"02F3", X"FF67", X"0010", X"FA80", X"F399", X"F44D", X"FE35", X"0034", X"FDC6", X"00BB", X"04FE", X"0AC5", X"0B64", X"06C2", X"00E7", X"FF77", X"FB3E", X"FE6F", X"FF2D", X"FED4", X"0174", X"0506", X"0505", X"04B9", X"011F", X"0194", X"024D", X"03B6", X"04A6", X"0211", X"020C", X"FC62", X"F3FA", X"F85C", X"FC83", X"FE2B", X"00C4", X"02D0", X"042F", X"0899", X"0C52", X"06BB", X"01C9", X"FF37", X"FC41", X"FD6E", X"FC5E", X"FCC6", X"0003", X"075A", X"0D73", X"09FF", X"05AA", X"041C", X"03FD", X"03BD", X"0346", X"02F8", X"031C", X"FC70", X"F3AE", X"F8B3", X"FDC4", X"0123", X"0090", X"02C0", X"0826", X"09EA", X"0B2F", X"06D1", X"0225", X"FD03", X"FC75", X"FAC6", X"FAEF", X"FA9F", X"FCF5", X"039C", X"0C37", X"081C", X"0636", X"04DF", X"047B", X"0450", X"03CF", X"018E", X"0098", X"FB99", X"F680", X"FDB8", X"FE4F", X"00A9", X"0222", X"0302", X"070C", X"0C59", X"0BC4", X"0535", X"FCC5", X"F7FE", X"FA00", X"F919", X"FB56", X"FB23", X"FA45", X"FBB8", X"05D8", X"05D4", X"023F", X"0227", X"02EF", X"044E", X"0174", X"FF4D", X"FC51", X"FAB6", X"F538", X"FCF9", X"FDE5", X"00D2", X"009C", X"0493", X"0749", X"0B4B", X"0B3E", X"0046", X"F868", X"F788", X"FC08", X"FBFB", X"FD6D", X"FB6E", X"F84C", X"F8A1", X"0299", X"0215", X"01DE", X"FF9F", X"013E", X"0134", X"FD47", X"FB1E", X"F71F", X"F505", X"FA0B", X"05D9", X"0606", X"03A4", X"0045", X"0044", X"05D4", X"08FB", X"0561", X"FD71", X"FAC8", X"FAEF", X"FB95", X"FE1E", X"FD1D", X"FA92", X"FA2D", X"FE36", X"01CC", X"0038", X"FF9F", X"037A", X"0262", X"FF5E", X"FD7A", X"FC28", X"F849", X"FA8F", X"FEF4", X"08C1", X"0924", X"0203", X"FCD0", X"0135", X"04B0", X"0A35", X"04A2", X"FEE7", X"FCD7", X"FE03", X"0044", X"FECC", X"FCF3", X"FBAD", X"FA96", X"FF33", X"02F7", X"010D", X"0047", X"00B4", X"0254", X"01B5", X"004A", X"FC2B", X"FC49", X"FE16", X"01F4", X"0788", X"08CD", X"02A3", X"FDB6", X"013B", X"02CA", X"0A2F", X"058D", X"0229", X"009B", X"FF21", X"FE3F", X"FD8C", X"FD19", X"FBAE", X"FD46", X"FFC9", X"0122", X"0113", X"0187", X"0140", X"01FE", X"FF4C", X"FFEE", X"FFE9", X"013A", X"014C", X"04FE", X"07B0", X"08E7", X"0400", X"00DF", X"0094", X"0186", X"092B", X"08FD", X"05DE", X"025A", X"FDBF", X"FC05", X"FE68", X"FD1B", X"FD24", X"FE88", X"0143", X"01B8", X"00AE", X"0306", X"014F", X"FFF0", X"FFD3", X"01AB", X"02FC", X"03F4", X"038D", X"0500", X"09A6", X"0A55", X"0460", X"FFC7", X"012C", X"01A0", X"096D", X"0AD9", X"04F1", X"0282", X"FDDD", X"FC87", X"FD4C", X"FD61", X"FAD2", X"FDA8", X"FF13", X"0079", X"0180", X"FF82", X"FF71", X"007C", X"008D", X"00F1", X"028B", X"0353", X"023C", X"03FE", X"09C0", X"0A33", X"0424", X"0302", X"00E8", X"0415", X"0896", X"0B3F", X"050E", X"0032", X"FE43", X"FCAA", X"FCBC", X"FD7D", X"FC53", X"FB2A", X"FECD", X"01F7", X"0050", X"0026", X"00D7", X"009D", X"01BA", X"0312", X"03D8", X"0462", X"0166", X"04DC", X"07A2", X"06E2", X"02C4", X"FFFF", X"023A", X"03C9", X"0433", X"0833", X"04DB", X"01A7", X"00C9", X"FD7A", X"00F2", X"FF5E", X"FB93", X"FCE2", X"FF42", X"008C", X"00EC", X"016E", X"024C", X"01BE", X"FFB1", X"00BF", X"0200", X"0060", X"0040", X"0193", X"07A3", X"0685", X"01B5", X"0006", X"FCC3", X"00DE", X"03E9", X"0789", X"060C", X"047C", X"02DC", X"012D", X"016E", X"FEA5", X"FFA4", X"FC83", X"FFA0", X"FF78", X"FF9A", X"0037", X"0043", X"0283", X"01D8", X"0136", X"027A", X"FFD9", X"009D", X"022A", X"0474", X"0635", X"FF7B", X"0047", X"00C7", X"0175", X"0259", X"04E6", X"049A", X"041C", X"01CA", X"0269", X"0184", X"0004", X"FE09", X"FD91", X"FC59", X"FEB0", X"FD57", X"0000", X"005E", X"023B", X"0298", X"01B5", X"0146", X"0006", X"005B", X"02D2", X"0424", X"0021", X"FF94", X"FEE9", X"018A", X"01B7", X"01FA", X"03DC", X"04AC", X"04DE", X"0445", X"0393", X"0156", X"01B7", X"FFC0", X"FCF2", X"FCF6", X"FC57", X"FE4D", X"FCD5", X"FF72", X"0253", X"0231", X"0482", X"0211", X"0297", X"01E0", X"FF5C", X"015B", X"FE40", X"FFA4", X"FFF5", X"01BC", X"0294", X"014F", X"0675", X"04AD", X"05EB", X"03BB", X"0138", X"00B0", X"015B", X"FF4F", X"FE7F", X"FD51", X"FC7D", X"FF27", X"FD19", X"FEDF", X"00D6", X"03A0", X"03BB", X"032B", X"02D0", X"FEE9", X"FF77", X"FFA4", X"0014", X"0069", X"FFA7", X"0028", X"00F8", X"00DD", X"047E", X"03A8", X"0403", X"03F7", X"0256", X"01B8", X"01A5", X"00DC", X"004F", X"0156", X"005F", X"FF1E", X"FDC2", X"FFCD", X"FD53", X"FED6", X"00CC", X"0383", X"0115", X"FEE9", X"01E8", X"0483", X"030C", X"FE93", X"0000", X"FFEA", X"FEBD", X"FDEE", X"017E", X"0440", X"02A1", X"01A2", X"03CA", X"03CA", X"0237", X"02E5", X"046F", X"040A", X"0383", X"01F1", X"0129", X"0174", X"01B5", X"00E8", X"0144", X"01E0", X"00E9", X"F812", X"FD73", X"026E", X"029B", X"0140", X"FF09", X"00B5", X"00E1", X"FE2B", X"FE2A", X"03C7", X"032E", X"0148", X"01D4", X"04BF", X"048F", X"020C", X"FF9D", X"028A", X"0531", X"0531", X"0708", X"05DF", X"04A6", X"04CA", X"022A", X"03A7", X"0400", X"0190", X"0037", X"FFBD", X"FFC6", X"003A", X"FF5E", X"00FE", X"FE78", X"0073", X"0079", X"027C", X"01BA", X"0232", X"0360", X"0278", X"0575", X"02EC", X"03B4", X"06B8", X"0608", X"0450", X"05CC", X"0731", X"0549", X"04C8", X"033A", X"04DF", X"037B", X"03D8", X"FFA6", X"0265", X"FF66", X"0009"),
        (X"FFD5", X"FFC4", X"FF5F", X"FFA6", X"010D", X"0086", X"0039", X"002D", X"FEE3", X"FEC9", X"01F8", X"FFCC", X"018A", X"009E", X"FED1", X"FF28", X"0042", X"FFCE", X"0080", X"001E", X"00B9", X"0058", X"FEFC", X"FFEB", X"0082", X"0066", X"0142", X"FFD9", X"FFD0", X"FEB7", X"FFFC", X"FF6B", X"0044", X"FFE3", X"04B0", X"061F", X"04A9", X"05E6", X"068A", X"09B6", X"08E5", X"0399", X"FF5F", X"0556", X"016F", X"03F2", X"05EA", X"0708", X"05AD", X"0353", X"02F2", X"0299", X"FFD7", X"0008", X"00A1", X"0039", X"0056", X"00B2", X"007F", X"00AD", X"0415", X"01E0", X"0628", X"0841", X"0941", X"0309", X"0750", X"075E", X"0823", X"066D", X"0751", X"0A6B", X"0B44", X"0A28", X"07F8", X"0729", X"07A6", X"070E", X"06B4", X"07BE", X"0538", X"010D", X"FEFC", X"FEE1", X"0107", X"0026", X"03B8", X"01CA", X"FF77", X"FE44", X"011E", X"0080", X"FD6B", X"FCCD", X"FD8F", X"FF06", X"FE83", X"010A", X"00A9", X"02DA", X"04B3", X"050D", X"04CC", X"052B", X"02BF", X"00DB", X"FDD4", X"0251", X"046D", X"0136", X"FEEA", X"01E3", X"0065", X"0036", X"0204", X"0285", X"FE54", X"FADC", X"FB3D", X"FA7B", X"FC21", X"FBA6", X"FC72", X"FBFE", X"FC0F", X"FE9F", X"000A", X"001B", X"FD1F", X"FF97", X"FE90", X"0115", X"0177", X"00A8", X"FE3D", X"FF3A", X"FC7D", X"FA2B", X"FDFC", X"020E", X"FFA7", X"00C8", X"00FF", X"FEEA", X"FA5A", X"F982", X"FB9A", X"FBFB", X"FED5", X"FEBE", X"FB7F", X"FC55", X"F9EE", X"FEAB", X"0037", X"FE99", X"FDC1", X"FF13", X"FFF0", X"FEE2", X"FCA2", X"FCB5", X"FAD8", X"F85B", X"F993", X"F522", X"FA53", X"0116", X"0105", X"003E", X"030C", X"00EA", X"FCE7", X"FC28", X"FE1E", X"FD50", X"00D5", X"FF5E", X"FF3B", X"FEC3", X"FDF4", X"FFDC", X"0121", X"002E", X"01FF", X"032E", X"03CE", X"FFC5", X"FEC9", X"FF93", X"FC7C", X"F9D1", X"F4FF", X"F0B6", X"F5F7", X"FC65", X"01E0", X"00B4", X"03DD", X"01DA", X"FDC3", X"FD6E", X"FEF2", X"FE80", X"FDF7", X"FE99", X"00C1", X"FF70", X"0008", X"01B2", X"022A", X"03B0", X"0308", X"06CB", X"04EA", X"01DD", X"0133", X"0067", X"FEC2", X"FDE3", X"F94F", X"F2B5", X"F327", X"FB99", X"026B", X"0416", X"026C", X"0360", X"FE8B", X"FF42", X"FF41", X"0041", X"0116", X"00DB", X"0073", X"FED9", X"FE8B", X"00BE", X"038E", X"0426", X"05A6", X"0593", X"03FE", X"0039", X"00AF", X"FDFE", X"FE31", X"FEA2", X"FAA8", X"F1E6", X"F308", X"FC53", X"0105", X"0551", X"02AA", X"0396", X"0013", X"FE6F", X"FFA3", X"FFFD", X"0177", X"FFF0", X"00F9", X"FCB5", X"FEA0", X"FFCC", X"02A3", X"04FA", X"059A", X"03BA", X"0215", X"FFCD", X"FE8D", X"FF24", X"FDC7", X"FF4D", X"FA50", X"F2BB", X"F9AB", X"02B4", X"022B", X"03AC", X"0606", X"03D6", X"007B", X"00A6", X"001F", X"0071", X"0104", X"FECA", X"FF38", X"FEB3", X"FCBA", X"FF35", X"04F5", X"0500", X"051C", X"01F2", X"0230", X"0038", X"0106", X"051B", X"0504", X"03A1", X"FA8C", X"F5D9", X"F9A6", X"0064", X"0173", X"0488", X"07CB", X"0445", X"0207", X"0008", X"0101", X"03A1", X"004D", X"FF9C", X"0035", X"FF51", X"FBD7", X"0033", X"02C3", X"0096", X"FF5A", X"0106", X"011B", X"FF8C", X"03AA", X"06D0", X"069A", X"0479", X"00B6", X"F339", X"F769", X"00C4", X"0131", X"0406", X"0804", X"043F", X"05E0", X"01FC", X"03B6", X"0452", X"0097", X"007F", X"FE43", X"FDE5", X"FBF1", X"F96E", X"FB58", X"FE25", X"FF83", X"0071", X"FF0C", X"014D", X"0134", X"0516", X"0929", X"090E", X"0A22", X"FAE4", X"FD80", X"0230", X"003F", X"034E", X"06AF", X"0451", X"05AA", X"0324", X"0343", X"00BC", X"011C", X"FEAE", X"FFF3", X"FE8E", X"FAF6", X"F8B8", X"F99E", X"FE19", X"FE37", X"FDFE", X"003C", X"0098", X"010C", X"053D", X"0836", X"0B51", X"0B6F", X"FFFE", X"FA2E", X"FD52", X"FDB8", X"00CA", X"04A2", X"02D5", X"02D4", X"0409", X"02BF", X"0213", X"01C3", X"01EE", X"0147", X"FE92", X"FEED", X"F9C7", X"FB48", X"FDF3", X"FC75", X"FE9B", X"021D", X"045B", X"039E", X"06B6", X"074C", X"086E", X"03F9", X"FDDC", X"F794", X"FDEA", X"FFCB", X"0121", X"FE87", X"FCE5", X"FFD2", X"031E", X"0329", X"03B2", X"029B", X"044F", X"02A9", X"00C0", X"FC9B", X"F9C6", X"FB32", X"FD15", X"FBB7", X"FFAF", X"01EF", X"045F", X"06A2", X"0526", X"0699", X"0660", X"00AA", X"FA9E", X"F97A", X"FC73", X"00F1", X"FE74", X"FC4A", X"F910", X"FE6B", X"017B", X"0143", X"0585", X"055A", X"05D6", X"0557", X"00E5", X"FB4E", X"F946", X"FACC", X"FC4E", X"FB1F", X"0014", X"02C0", X"019A", X"010F", X"0139", X"0204", X"FEEB", X"FD83", X"F856", X"F99E", X"FD44", X"FEC1", X"0051", X"FACA", X"F688", X"FB7D", X"FE3F", X"0079", X"FE58", X"01AB", X"0434", X"052F", X"012D", X"FCAB", X"FE56", X"FD2D", X"FBF2", X"FC5C", X"FD84", X"FCB4", X"FD27", X"FF75", X"000C", X"0068", X"FE57", X"FB6D", X"FFFB", X"FDD1", X"00C9", X"01E0", X"FFFA", X"FCF3", X"F4D5", X"FA7C", X"FC2D", X"FC98", X"FDC8", X"FEF2", X"01E5", X"03FB", X"0316", X"FFE2", X"0132", X"FD32", X"FB23", X"FA79", X"FD06", X"FD2E", X"FDAD", X"FD5B", X"FE19", X"FE58", X"F9EB", X"F8ED", X"FFC5", X"00A2", X"FC6B", X"0025", X"0471", X"FEF5", X"F7E0", X"FB76", X"F9EE", X"FB37", X"FD8A", X"FC25", X"00A3", X"02C4", X"06F7", X"0768", X"030B", X"FF7F", X"FC31", X"F9BE", X"FC0E", X"FCF8", X"FB97", X"FC7F", X"FCB5", X"FAEF", X"F9BA", X"FB31", X"FED5", X"FF05", X"0209", X"010B", X"0286", X"FBFA", X"F9B7", X"F794", X"FC8D", X"FA52", X"FBCB", X"FB93", X"FD6A", X"02E4", X"0737", X"07BE", X"03E9", X"0395", X"FF19", X"FBA3", X"FABA", X"F900", X"FA8D", X"F9EF", X"FA54", X"F7B4", X"F8F2", X"FE49", X"FF1F", X"0026", X"0017", X"016B", X"00A2", X"FB8C", X"FAF5", X"FBA5", X"FB3A", X"FD23", X"FCA5", X"FDBE", X"FFF1", X"0218", X"0377", X"037D", X"0213", X"0482", X"00BF", X"FF4E", X"F97C", X"FA1F", X"F8CF", X"F8E5", X"FB2B", X"F54C", X"F83A", X"FE96", X"0066", X"02DC", X"FFE0", X"00D2", X"0087", X"FB36", X"F70E", X"F9CF", X"FFAC", X"FE42", X"FFA1", X"007C", X"0010", X"FE1A", X"0106", X"FF9B", X"00B0", X"01E8", X"029A", X"FED0", X"FC2E", X"F847", X"F7F1", X"F764", X"F65A", X"F610", X"F82C", X"FBC1", X"FDA4", X"0196", X"FFEF", X"0126", X"FFD1", X"FADA", X"F808", X"FCCC", X"0042", X"0037", X"01F1", X"0086", X"012C", X"FF88", X"FDF2", X"0155", X"0251", X"0317", X"0414", X"FDF9", X"FB78", X"F6BC", X"F3F4", X"F2DE", X"F492", X"FA29", X"F61B", X"FB4B", X"FC8B", X"01A2", X"00DB", X"FFCC", X"008B", X"FF69", X"0087", X"02E1", X"05C5", X"033F", X"0176", X"007B", X"FDFD", X"FE08", X"FC66", X"FCDF", X"FE37", X"FDE5", X"0093", X"FEC1", X"FDD8", X"F9C4", X"F72B", X"F826", X"FAE7", X"F91A", X"F8F3", X"FBBD", X"FC3D", X"01AE", X"FFC6", X"FEFF", X"0057", X"FDF7", X"026C", X"068B", X"0406", X"027E", X"0184", X"007B", X"FD78", X"FD24", X"0081", X"00D4", X"00DE", X"017C", X"0431", X"03C0", X"0504", X"0340", X"0514", X"02E6", X"0455", X"004D", X"FBCE", X"FEB8", X"0051", X"FED1", X"FF8D", X"FF3B", X"010A", X"00C0", X"FE3A", X"FEDF", X"02D9", X"00AA", X"005C", X"00CF", X"0310", X"0231", X"02E5", X"0167", X"0575", X"0717", X"04C8", X"06BC", X"0702", X"0A2C", X"0B5F", X"0618", X"0514", X"02CB", X"FF0D", X"015C", X"0007", X"0020", X"FF4B", X"FE70", X"FEB5", X"FF46", X"0034", X"0139", X"0011", X"026F", X"0460", X"03BA", X"036C", X"0544", X"03F1", X"03CE", X"09C7", X"03ED", X"0324", X"059F", X"09F7", X"07D2", X"0525", X"0337", X"02BB", X"0187", X"032A", X"FFF9", X"FFAF", X"007C", X"00A4"),
        (X"FF8A", X"0079", X"000C", X"0071", X"FF5F", X"FFD1", X"FF0F", X"FE8B", X"00D4", X"00DB", X"FFA2", X"FFF4", X"00CE", X"FEC9", X"FFD6", X"00D5", X"FF64", X"000C", X"0066", X"FFC5", X"FF0E", X"FF20", X"FF8B", X"00B5", X"FFA0", X"FF78", X"0014", X"FF90", X"0047", X"00AE", X"0062", X"00F2", X"0162", X"0127", X"00B1", X"0261", X"0291", X"02DB", X"01E8", X"0262", X"0090", X"FF74", X"FEA1", X"FDDE", X"FBCF", X"FE78", X"039A", X"0526", X"03D1", X"02EF", X"03E7", X"FFB1", X"FF09", X"FF06", X"00F8", X"005B", X"0027", X"FEC0", X"00FC", X"FC4B", X"FE3A", X"0171", X"0226", X"0130", X"04DF", X"05DA", X"0608", X"02F8", X"0202", X"005E", X"0114", X"00B8", X"FF85", X"04C4", X"0533", X"07AE", X"084C", X"071C", X"06F4", X"0548", X"0104", X"007A", X"FF8A", X"0055", X"FF48", X"FFED", X"FDF8", X"FDD3", X"0235", X"018F", X"03F5", X"03E7", X"03B2", X"02B1", X"0317", X"0065", X"FCBA", X"FD08", X"FDA2", X"FCE6", X"FA3A", X"FE30", X"0151", X"05EB", X"0587", X"07B7", X"07AB", X"0525", X"055A", X"031A", X"0079", X"FFD7", X"0122", X"FFBA", X"FD69", X"0031", X"02C9", X"02BA", X"01C7", X"023A", X"FFE5", X"00A8", X"FEF7", X"FD0E", X"FAED", X"F9EA", X"F868", X"F61D", X"F8A8", X"FC72", X"FF86", X"FE3F", X"0039", X"0387", X"0458", X"09DC", X"0948", X"02B2", X"FC30", X"FEE5", X"FE76", X"00EE", X"FD64", X"01FD", X"0045", X"0369", X"0329", X"0389", X"0295", X"026E", X"02BA", X"0055", X"FFC6", X"FD90", X"FB44", X"F84A", X"F969", X"FA33", X"FC3B", X"FEAE", X"FEF4", X"00A6", X"02D5", X"0608", X"0628", X"01DB", X"0122", X"0347", X"00F6", X"FF01", X"0032", X"FEBE", X"03E1", X"0189", X"0448", X"04D0", X"03B7", X"02B3", X"0154", X"0177", X"FFC9", X"FF6C", X"FE37", X"FBBE", X"F941", X"FBA5", X"FBAB", X"FD54", X"FE6C", X"FD53", X"FE0E", X"043B", X"05FC", X"03FB", X"0608", X"03B7", X"FFEE", X"FD03", X"000A", X"FEF1", X"FE68", X"008A", X"01BA", X"02F6", X"0288", X"026E", X"009C", X"038A", X"003C", X"FFAE", X"0001", X"FECE", X"FC33", X"FB6F", X"FB39", X"FD31", X"FE94", X"FE50", X"FC74", X"0043", X"04CC", X"0715", X"0209", X"01EB", X"FC3F", X"FDCB", X"0257", X"FE86", X"FE93", X"00ED", X"FFB9", X"FFFA", X"0156", X"01D9", X"02F1", X"036E", X"011F", X"0289", X"0116", X"FCF4", X"F9EA", X"F7F5", X"F9D0", X"FCD2", X"FE71", X"FD92", X"FC59", X"FFFB", X"06D5", X"07EC", X"01A7", X"FF74", X"0067", X"040D", X"FFAA", X"FE0D", X"00C3", X"00AC", X"0232", X"0267", X"04CD", X"02A4", X"03DB", X"043D", X"03CF", X"0442", X"050A", X"FF2C", X"FB8F", X"F8C0", X"F86B", X"F904", X"FB71", X"FD25", X"FD2A", X"000B", X"0875", X"0AAE", X"0413", X"01EE", X"FF77", X"02FE", X"FDE2", X"0160", X"0261", X"0357", X"0490", X"0334", X"040B", X"046D", X"0468", X"04B2", X"0784", X"0919", X"05AE", X"00B8", X"FDF8", X"FBD2", X"F934", X"FA5A", X"FA86", X"FB02", X"F82C", X"FDBF", X"07AC", X"0D6C", X"06A8", X"FD69", X"FF18", X"FDC9", X"0204", X"04D4", X"0763", X"0759", X"0671", X"050C", X"042D", X"03E9", X"03DA", X"02BA", X"06DC", X"06EB", X"00F0", X"FFAC", X"01CC", X"0217", X"FDF6", X"FC3C", X"FB02", X"F913", X"F785", X"F766", X"FF4C", X"06BC", X"0480", X"FE00", X"004C", X"00D5", X"04E0", X"0875", X"08D0", X"09B6", X"06BF", X"061A", X"0373", X"013C", X"005F", X"0260", X"03F7", X"027F", X"010F", X"FD18", X"004D", X"01BF", X"0186", X"FEB3", X"FE20", X"FA2C", X"F82A", X"F68D", X"F558", X"FDAA", X"FD2D", X"FB16", X"FDFB", X"FF87", X"0172", X"0512", X"08FD", X"066D", X"0496", X"0283", X"002B", X"FF3D", X"00C4", X"0116", X"02D1", X"0045", X"FD83", X"FE91", X"01E3", X"026B", X"01CA", X"00FF", X"0064", X"FE7F", X"FD3B", X"FB8A", X"FAE6", X"FDC3", X"FAC1", X"FD4E", X"0168", X"01CA", X"00C0", X"05F9", X"04FF", X"FF9C", X"FFF1", X"FCC9", X"FE5E", X"FE77", X"FF90", X"00A4", X"0161", X"FE15", X"FE67", X"FF5B", X"030F", X"0070", X"FF55", X"000F", X"003A", X"FF0E", X"004D", X"003D", X"00F6", X"00FD", X"FA2D", X"FE2D", X"00E4", X"FF52", X"FE57", X"0177", X"FC9B", X"F9E5", X"FEB5", X"FBA4", X"FCAB", X"FD7C", X"FFBE", X"0206", X"00CF", X"FD5C", X"FFF4", X"0293", X"03C1", X"03C6", X"0158", X"00A0", X"014B", X"007D", X"01FE", X"FFD4", X"021D", X"021E", X"FD7F", X"FD43", X"005C", X"FF18", X"FC40", X"FF04", X"FB2A", X"F79C", X"FCBC", X"FC52", X"FBD3", X"FA53", X"FC8A", X"FF08", X"FECB", X"0174", X"05CF", X"05B4", X"043B", X"03A6", X"02C5", X"04B2", X"021D", X"007E", X"00D7", X"023A", X"031D", X"0113", X"FC6F", X"FCB1", X"0004", X"FEDE", X"FE69", X"FFAD", X"FDEF", X"FC9F", X"FF91", X"FEDE", X"FBC2", X"FA4F", X"FBED", X"FCA6", X"FDEA", X"037E", X"08BF", X"0767", X"0234", X"037B", X"031B", X"02E8", X"0545", X"024B", X"0220", X"007B", X"0084", X"FE28", X"FB15", X"FC18", X"FE5B", X"FE66", X"00E2", X"00E2", X"FEC0", X"FEAD", X"00EB", X"FFC5", X"FDB2", X"FA8F", X"F98F", X"FDA8", X"035E", X"0888", X"0A40", X"04BD", X"0429", X"0323", X"0164", X"045C", X"02BC", X"02B7", X"FFC8", X"FF7F", X"FCDD", X"FBF7", X"FD4B", X"FC7D", X"005B", X"FD7D", X"00D5", X"00BC", X"0011", X"FEE0", X"0144", X"FE4A", X"FDBD", X"FAFB", X"F959", X"FC31", X"0380", X"0740", X"0513", X"01DF", X"02B7", X"02B8", X"032C", X"0342", X"02EF", X"014D", X"FE4B", X"FE74", X"0029", X"FBD2", X"FB1C", X"FCF7", X"FEF5", X"FD2F", X"01EC", X"FFA4", X"FFE6", X"FF72", X"FDC0", X"FC17", X"FC31", X"FAE3", X"FA59", X"FE55", X"0259", X"051F", X"04AF", X"01E7", X"03FB", X"0305", X"03F8", X"0209", X"014A", X"FF3F", X"FF41", X"FEDD", X"FF5E", X"FFF8", X"FB2F", X"FF73", X"00A8", X"FE9B", X"FA99", X"0010", X"029D", X"FF36", X"FCAB", X"FD09", X"FE7E", X"FDA9", X"FDAC", X"FED5", X"02C6", X"0174", X"01A9", X"0346", X"0418", X"03F4", X"01AC", X"033B", X"0220", X"0179", X"0248", X"0189", X"0306", X"0192", X"FC6B", X"0066", X"0084", X"FF7E", X"FA2B", X"FEFC", X"0240", X"FDCA", X"FA2B", X"FB68", X"FD1F", X"FD0A", X"FD7A", X"FDDB", X"00AC", X"FFB9", X"FE22", X"014D", X"0313", X"02A0", X"01D0", X"036F", X"0330", X"0247", X"00F7", X"028A", X"048C", X"0306", X"0029", X"FFC1", X"0099", X"0068", X"FB9B", X"0003", X"00C7", X"FFA2", X"FC8C", X"FBA7", X"FBAF", X"FD93", X"FE60", X"FEA4", X"FB30", X"FBF5", X"FEE9", X"FFA1", X"00DD", X"FFE5", X"00C6", X"03E5", X"0484", X"0537", X"03DA", X"0344", X"02E5", X"03D7", X"00BD", X"00BB", X"FFC2", X"FF17", X"FE7C", X"FAE5", X"FAF0", X"FFB4", X"FF99", X"0115", X"0023", X"00F4", X"FFD5", X"FE4F", X"FD1D", X"FDBE", X"FFA6", X"FF58", X"FF95", X"0153", X"0472", X"05FF", X"0581", X"0426", X"0730", X"0599", X"FFD5", X"FBB2", X"FE21", X"00B6", X"0109", X"008C", X"FF33", X"FF10", X"FFA7", X"0138", X"0016", X"0019", X"009C", X"021A", X"FFA0", X"0031", X"024B", X"01CA", X"0241", X"02DF", X"05B0", X"0686", X"056A", X"05DF", X"05EC", X"040F", X"05FE", X"04F7", X"04A4", X"FF9D", X"FE57", X"00F4", X"00D6", X"FE47", X"0199", X"011B", X"045C", X"0519", X"07A8", X"064E", X"05BA", X"05B3", X"075B", X"083C", X"09AD", X"0772", X"06AE", X"07B7", X"0518", X"04D5", X"0536", X"05BB", X"0582", X"0393", X"0030", X"FF67", X"0049", X"0202", X"001A", X"0097", X"0006", X"00CA", X"FFD3", X"FECC", X"005D", X"00AC", X"0137", X"FEAE", X"0062", X"02A6", X"0435", X"040E", X"035C", X"03C1", X"03C6", X"02D2", X"0266", X"026C", X"00F8", X"01E0", X"FFD5", X"0159", X"01FF", X"FFCE", X"FFE4", X"FF90", X"003E", X"FF80"),
        (X"00E4", X"0098", X"FFA4", X"01AB", X"FF7E", X"0107", X"00D6", X"FF9F", X"011A", X"FFD8", X"00B9", X"009D", X"FDEC", X"FCEE", X"0108", X"FF12", X"FF89", X"0129", X"FFC0", X"FF0D", X"0165", X"008F", X"00FD", X"0103", X"FF9D", X"FF9F", X"00D0", X"FF67", X"FFC0", X"0065", X"009F", X"FF31", X"00C3", X"FDDD", X"FC06", X"FBD7", X"FD02", X"FD0C", X"FC78", X"FEA5", X"0056", X"FE4F", X"FD12", X"FC31", X"03D6", X"00A4", X"FAFC", X"FCFE", X"FB30", X"FDB4", X"FEAE", X"FE9F", X"0182", X"FFD4", X"00D8", X"0006", X"0045", X"003C", X"0021", X"0227", X"FF75", X"FCA9", X"FCD9", X"FBD0", X"FDEC", X"FDAF", X"FA27", X"FA12", X"FB7C", X"FB26", X"FB8F", X"FCC9", X"FE3C", X"FEF6", X"FDF8", X"FBEA", X"F9A6", X"F748", X"F7F6", X"FAC2", X"FDDA", X"00F9", X"FF9E", X"FFBC", X"0071", X"00E1", X"FFA0", X"007A", X"01F4", X"FFC0", X"FD0B", X"FDF9", X"FD42", X"FDA4", X"FF0C", X"0056", X"036C", X"0246", X"017B", X"0093", X"0005", X"FEAC", X"FDFF", X"FDB7", X"FDB8", X"FB8F", X"F8CC", X"F990", X"FC77", X"FF80", X"0011", X"008D", X"006F", X"011B", X"FEB9", X"00D1", X"0097", X"003A", X"FFE2", X"006C", X"00F3", X"00F6", X"0182", X"0649", X"06A7", X"0654", X"0583", X"06B8", X"00B7", X"0030", X"006A", X"FC97", X"F934", X"F962", X"F87C", X"FC44", X"0154", X"03AD", X"0241", X"FE2B", X"FFFF", X"FEEA", X"FDA8", X"FFD1", X"FFF1", X"0005", X"0225", X"0415", X"04BF", X"05E7", X"0588", X"0717", X"0485", X"048C", X"0416", X"0395", X"0499", X"03C4", X"025C", X"FDBF", X"FC0C", X"FC52", X"FEC2", X"FFDC", X"0114", X"04AB", X"0242", X"FE12", X"002E", X"000E", X"01DF", X"0100", X"0206", X"0626", X"04B7", X"064D", X"08A1", X"0527", X"061A", X"0276", X"026B", X"0147", X"00A8", X"FFB6", X"019D", X"011B", X"0094", X"FF8C", X"FDFF", X"FF99", X"0312", X"040E", X"05F7", X"079A", X"02C1", X"FE16", X"FF9B", X"0259", X"019A", X"0336", X"04EB", X"0746", X"0898", X"0827", X"0A04", X"0305", X"0240", X"0149", X"FF46", X"FE90", X"FE4A", X"FF54", X"00E5", X"023E", X"0334", X"FF0E", X"FE87", X"0073", X"01D9", X"051F", X"0690", X"0827", X"03A1", X"FF4E", X"02C5", X"024D", X"0471", X"05E1", X"03C0", X"059D", X"075E", X"07D8", X"0585", X"031C", X"00F7", X"02B4", X"FF78", X"002D", X"0133", X"029A", X"052D", X"03CA", X"0354", X"02F6", X"039F", X"01EA", X"0203", X"0535", X"053D", X"05C2", X"063F", X"029A", X"02CC", X"01B1", X"04E8", X"05EA", X"0649", X"0851", X"077E", X"0553", X"0320", X"01FB", X"0161", X"0188", X"01AD", X"0088", X"FFC4", X"018F", X"0526", X"054C", X"052C", X"052A", X"060D", X"04E2", X"03B5", X"06A6", X"0815", X"0A97", X"09EE", X"0482", X"022E", X"011E", X"0562", X"0746", X"05CE", X"07B7", X"0889", X"04A2", X"008E", X"01B9", X"FEFC", X"FFE4", X"FE65", X"FD1F", X"FDDD", X"FE4C", X"0383", X"056B", X"0514", X"0336", X"067F", X"05B2", X"0615", X"0BEB", X"0DC3", X"0D28", X"0914", X"FFEF", X"FFF6", X"04A9", X"05D0", X"0759", X"07BB", X"0675", X"046E", X"0223", X"FCE9", X"FB0A", X"FCB0", X"FC3A", X"FBDB", X"FC9E", X"FC1C", X"FDBB", X"FECE", X"01DA", X"0272", X"0321", X"024B", X"FD8E", X"011F", X"0704", X"0B18", X"0CB6", X"0798", X"FD9E", X"FF62", X"02AD", X"0408", X"0569", X"042B", X"058C", X"01D6", X"FDDB", X"FCCA", X"FAE9", X"FB20", X"FBC6", X"FBFD", X"FBB4", X"FBC4", X"FBED", X"FD30", X"0003", X"011D", X"FF6D", X"FBC2", X"F521", X"F7B0", X"FC09", X"01FB", X"057A", X"0656", X"01A4", X"001F", X"0212", X"04CF", X"03DC", X"01D1", X"03E5", X"0254", X"000B", X"FAE3", X"FB43", X"FCB2", X"FFAF", X"011A", X"FF98", X"FC3D", X"FB8B", X"FBDE", X"FDF4", X"FD76", X"FBBD", X"F789", X"F456", X"F6F5", X"FE9D", X"027F", X"05FF", X"07D6", X"02DA", X"0039", X"00AE", X"0416", X"029C", X"0178", X"0452", X"02FB", X"FFC0", X"FCBF", X"FBD6", X"FE33", X"00BE", X"010D", X"FEE5", X"FBAA", X"F977", X"FB16", X"FD24", X"FFA2", X"FD7A", X"FB6E", X"FA7F", X"FCAF", X"010F", X"0638", X"05FF", X"0836", X"03AE", X"0144", X"FFD3", X"005F", X"044A", X"0411", X"0701", X"0692", X"FE95", X"FCD1", X"FE29", X"FE7C", X"FF09", X"FFE1", X"FE47", X"FB8E", X"FB0E", X"FB00", X"FFB7", X"01D2", X"0355", X"00E6", X"0142", X"03D9", X"0584", X"08D3", X"0703", X"07FB", X"010C", X"FF95", X"FFD2", X"00E4", X"0687", X"0581", X"0A82", X"09E3", X"0036", X"FCE0", X"FF38", X"FD2F", X"FDF3", X"0122", X"FDF0", X"FB6E", X"FB9F", X"FE98", X"02DC", X"0669", X"050D", X"04EC", X"0631", X"0692", X"0914", X"0B7E", X"09A8", X"06EC", X"03BA", X"FF36", X"FF19", X"023F", X"0809", X"06CC", X"0D0D", X"0B82", X"06DA", X"FEDF", X"FE3F", X"FB3B", X"FBFA", X"FD17", X"FE0C", X"FAD9", X"FD56", X"00C4", X"0430", X"062D", X"06E5", X"05F2", X"0550", X"0762", X"072A", X"0C11", X"0A07", X"0602", X"057A", X"FFF5", X"012B", X"0362", X"03E8", X"0960", X"0B97", X"0D6A", X"089A", X"0393", X"FDC8", X"FC13", X"FCEE", X"FCFD", X"FE6A", X"004D", X"FF47", X"03A2", X"03FE", X"02F3", X"031E", X"0334", X"046F", X"08FF", X"0911", X"0BA2", X"0748", X"FF37", X"00E3", X"0066", X"02D8", X"0407", X"0340", X"062C", X"07E7", X"0999", X"06D6", X"047A", X"0047", X"FDEC", X"FBB9", X"FF31", X"FFF2", X"0145", X"02AA", X"0170", X"0143", X"014F", X"01BF", X"02A8", X"0455", X"086E", X"08B1", X"08F9", X"0507", X"0170", X"FD87", X"FEDF", X"0266", X"044D", X"0703", X"07E3", X"0905", X"0816", X"0463", X"0345", X"FF3F", X"FE48", X"FE62", X"FDB9", X"FF1E", X"0046", X"0126", X"0129", X"FFE3", X"014C", X"01D2", X"032A", X"0351", X"05E9", X"062C", X"080C", X"0575", X"FE46", X"FF70", X"FFCA", X"FF27", X"03D9", X"035A", X"0859", X"069B", X"0484", X"01DE", X"FF88", X"FF08", X"FD65", X"FF69", X"FF09", X"FEA1", X"FF63", X"FEF8", X"FF7A", X"FFC6", X"FF0A", X"0381", X"035C", X"020F", X"06D0", X"0598", X"0006", X"0473", X"01AD", X"0133", X"FFAF", X"FFE9", X"FF9D", X"029F", X"0590", X"01B8", X"011D", X"03C9", X"0056", X"00A3", X"014B", X"0093", X"01AD", X"010C", X"005C", X"FFF5", X"FEF1", X"FE9C", X"FF61", X"025F", X"044C", X"048B", X"04DE", X"0353", X"007E", X"0143", X"011F", X"FFDE", X"FE6F", X"FF8B", X"0382", X"04D2", X"03BA", X"0002", X"FEFE", X"0156", X"020E", X"028E", X"0350", X"0334", X"0117", X"01AF", X"01AB", X"0262", X"FF41", X"FF73", X"0068", X"02C7", X"04B6", X"0547", X"031C", X"007D", X"00EA", X"013F", X"FF97", X"0046", X"FF32", X"FE6B", X"023E", X"045B", X"027D", X"FD88", X"00A5", X"00C3", X"0147", X"0241", X"0213", X"0204", X"049A", X"066C", X"06CC", X"0353", X"0172", X"00D0", X"FF8A", X"0190", X"0108", X"FE91", X"FE02", X"FCD2", X"0209", X"01CA", X"0195", X"0016", X"009F", X"00CF", X"FDD7", X"FC9E", X"FDA6", X"FCEC", X"FF46", X"00AA", X"0010", X"0253", X"00FD", X"0060", X"02E8", X"0341", X"0067", X"032A", X"0315", X"01E3", X"FFB9", X"0199", X"FEBE", X"FF4B", X"0147", X"FFE3", X"FE50", X"030B", X"022F", X"FFA6", X"00C1", X"FFBD", X"FF3B", X"FE01", X"FD02", X"FA96", X"F84B", X"FBF7", X"0056", X"FE75", X"FE1E", X"FE48", X"FF70", X"0142", X"FD8A", X"00D6", X"0054", X"0161", X"FFA4", X"00A9", X"FE6C", X"FEC0", X"0163", X"FF64", X"FF1F", X"0339", X"FFDC", X"FFA6", X"01E1", X"008C", X"FFCE", X"0101", X"013C", X"04E6", X"01BE", X"FFDF", X"012D", X"032D", X"02EF", X"018E", X"FF9D", X"0608", X"FF62", X"0047", X"0291", X"047E", X"00C8", X"0030", X"0039", X"007C", X"FF63", X"00B3", X"FF38", X"FECC", X"00A7", X"001F"),
        (X"0043", X"FFA9", X"FFA8", X"FEF1", X"0088", X"FF15", X"FFB8", X"0093", X"FF45", X"FFFA", X"0093", X"FF21", X"FFEB", X"FFFA", X"00E4", X"FFC4", X"FFCB", X"0000", X"009A", X"0050", X"004B", X"016C", X"FF47", X"00B6", X"FE61", X"0106", X"0019", X"0034", X"FE33", X"FF23", X"0114", X"FF91", X"FF95", X"FE93", X"FD7D", X"FCB5", X"FE13", X"FD00", X"FBFF", X"FB2D", X"FB45", X"FC99", X"00F7", X"01D8", X"0350", X"FEC9", X"FCA8", X"FDCD", X"FC0E", X"FE84", X"FECE", X"FF09", X"FFDF", X"FFCE", X"0013", X"FE4E", X"008D", X"002C", X"FFE7", X"FFF3", X"011C", X"FF56", X"FD2B", X"FBF7", X"FCC4", X"FFDD", X"FCF2", X"FE2E", X"0024", X"FFB8", X"001D", X"0088", X"0389", X"003E", X"FC97", X"FB79", X"FD01", X"FC97", X"FDD0", X"FFFE", X"017C", X"0307", X"0066", X"FFBC", X"007C", X"0179", X"021B", X"010C", X"FCA2", X"0152", X"FFF7", X"FF5B", X"FEC1", X"006E", X"01FC", X"0283", X"0621", X"054A", X"05B9", X"040D", X"022D", X"FF28", X"FC32", X"FB08", X"FCAD", X"F7A4", X"F6A3", X"F958", X"FA98", X"FD62", X"FF09", X"00DD", X"00B5", X"FF70", X"0266", X"0242", X"00CC", X"027F", X"04FD", X"02DD", X"0325", X"0331", X"0572", X"0447", X"0548", X"06DC", X"0396", X"037E", X"012B", X"FFB0", X"FE32", X"FFAC", X"FD23", X"F99D", X"FA4B", X"FA91", X"FA76", X"F90F", X"FBAE", X"FC93", X"0021", X"FEB7", X"01C6", X"0454", X"0364", X"04D8", X"06B3", X"05D4", X"0522", X"03F6", X"0567", X"0236", X"0159", X"01B9", X"00B7", X"0175", X"0104", X"FDA4", X"FEDB", X"FEBE", X"FCC9", X"FB39", X"FC94", X"F9E3", X"FD3D", X"F6BF", X"FAB9", X"FD17", X"0141", X"0146", X"0168", X"0681", X"051D", X"0657", X"0680", X"03D2", X"0529", X"03DD", X"0480", X"028E", X"011B", X"016A", X"FFA3", X"0015", X"FE33", X"FFC4", X"00FC", X"0065", X"0153", X"FFB4", X"FBC8", X"FA51", X"F8CF", X"F658", X"FD6D", X"FD25", X"FE6B", X"0292", X"009A", X"05DC", X"088B", X"0836", X"065F", X"01E8", X"005E", X"01BF", X"017C", X"017C", X"020F", X"000E", X"FF11", X"FD57", X"FF63", X"007B", X"0102", X"02A8", X"0289", X"019D", X"0011", X"FA0E", X"F627", X"F54A", X"FD3A", X"FF1E", X"FD16", X"0536", X"0436", X"058C", X"0790", X"035B", X"0234", X"0036", X"FF4D", X"FFBF", X"0170", X"037E", X"04D9", X"0348", X"0241", X"0179", X"013E", X"029F", X"0383", X"049A", X"0419", X"0014", X"012D", X"F71A", X"F5A6", X"F6EA", X"FBD6", X"FEF5", X"00CD", X"03D8", X"03E7", X"05D9", X"06D6", X"0234", X"00AD", X"024F", X"000D", X"FEFC", X"FF0B", X"010F", X"024A", X"06EF", X"0651", X"0638", X"0367", X"0354", X"0368", X"042A", X"01AA", X"000F", X"FCC0", X"F7F1", X"F500", X"F98C", X"FBF9", X"0100", X"0175", X"0444", X"071F", X"0781", X"0392", X"01B9", X"00D1", X"FE4B", X"FAE6", X"FBF3", X"FCBC", X"FDE4", X"0014", X"07AD", X"098E", X"0514", X"0459", X"0367", X"02B8", X"0366", X"0189", X"00F5", X"FB31", X"F7DA", X"F78A", X"FE50", X"FF24", X"00D3", X"003E", X"0477", X"085C", X"08C3", X"02C3", X"FD73", X"FDBD", X"FDC3", X"FB7E", X"FB3A", X"FB4E", X"FB3B", X"FC23", X"0328", X"05ED", X"0277", X"0266", X"000D", X"02F4", X"FFE9", X"FECB", X"FC00", X"FAB3", X"F852", X"F6B1", X"FF22", X"FDCE", X"00DF", X"007A", X"0556", X"053D", X"0362", X"027C", X"FE22", X"FAAC", X"FE24", X"FDC4", X"FC09", X"FA65", X"F6C2", X"F75C", X"FC02", X"0363", X"0234", X"FE9B", X"FFCE", X"FFED", X"FD16", X"FAF2", X"F7D5", X"F6DE", X"F6B0", X"F843", X"04E9", X"03D3", X"035C", X"0028", X"036B", X"0759", X"02D2", X"FEFD", X"FAB3", X"FB89", X"FB50", X"FB67", X"FB55", X"F826", X"F5A2", X"F44C", X"FC42", X"FFB5", X"FF2D", X"FEE9", X"FF1C", X"FFFF", X"FE5D", X"F9CA", X"F954", X"F5BD", X"F705", X"FBE5", X"05F2", X"04F3", X"01B6", X"FE8D", X"0174", X"0386", X"01D5", X"FDB4", X"F6D2", X"F6E2", X"F9CD", X"FA05", X"F843", X"F89F", X"F505", X"F818", X"FBC9", X"004B", X"FFAC", X"FE99", X"FFF4", X"0238", X"0123", X"FE5B", X"FBB3", X"FB7A", X"FBA0", X"FD65", X"054F", X"08F5", X"0223", X"FF96", X"0006", X"053E", X"FFB2", X"FAFC", X"F6B1", X"F7A5", X"F7A0", X"F95B", X"F8D5", X"F886", X"F9DE", X"FB69", X"01B9", X"0174", X"00AC", X"FED6", X"0052", X"01F3", X"0202", X"0249", X"FFD0", X"005B", X"0079", X"031B", X"047E", X"06C8", X"04A1", X"0252", X"0107", X"0553", X"0119", X"FACD", X"F6E9", X"F88B", X"F842", X"F935", X"FBB9", X"FB06", X"FCBE", X"FEDB", X"02CE", X"0150", X"FE1C", X"FF5A", X"FF7B", X"007F", X"00AF", X"0190", X"0402", X"0449", X"005E", X"03A5", X"0546", X"0829", X"04DA", X"00EE", X"0061", X"0562", X"0216", X"FC96", X"F871", X"F6E8", X"FA11", X"FA8B", X"FBB4", X"FE7C", X"FDAA", X"0021", X"0407", X"FF4F", X"00D4", X"FEC2", X"FEBE", X"FF7A", X"FFF5", X"0128", X"0163", X"0450", X"03B6", X"0379", X"0987", X"09B0", X"04C3", X"03D6", X"0116", X"0449", X"052E", X"FFE3", X"FB57", X"FBCD", X"FC17", X"FD46", X"FC7C", X"FBC3", X"FE07", X"0172", X"00B2", X"0262", X"01CF", X"FFAF", X"00F2", X"009F", X"0041", X"01E0", X"0385", X"03A9", X"0241", X"002E", X"0657", X"0750", X"047D", X"FF3A", X"01E5", X"046D", X"067A", X"00B0", X"FBD2", X"FCE0", X"FE64", X"FEC7", X"008F", X"FFBD", X"00A1", X"02CB", X"0108", X"0164", X"FFAE", X"00C4", X"0206", X"00E4", X"00E1", X"00D9", X"01EB", X"0229", X"0120", X"0171", X"07A7", X"07B6", X"025F", X"000F", X"FD93", X"01A8", X"0719", X"021E", X"FFF9", X"00B0", X"00CC", X"00B1", X"01FB", X"00DC", X"014D", X"FF93", X"FFF3", X"0102", X"0093", X"002D", X"0145", X"02C3", X"0132", X"014F", X"00C9", X"FF9D", X"FF7D", X"03B5", X"053E", X"0415", X"0149", X"0148", X"FFFE", X"0257", X"0711", X"05A9", X"042D", X"025D", X"00E5", X"03CF", X"005A", X"019B", X"FEFF", X"FEBE", X"FE4F", X"FF91", X"0245", X"01B7", X"012E", X"0137", X"0134", X"FFBF", X"FDD1", X"FD00", X"0152", X"02CA", X"0487", X"0383", X"0027", X"FF9C", X"FEFA", X"0393", X"04D9", X"04F4", X"06B6", X"0632", X"0350", X"029B", X"021A", X"0087", X"FFE3", X"FF8E", X"FC77", X"007E", X"01A3", X"0015", X"014B", X"0223", X"0186", X"FF08", X"FD89", X"FBF6", X"FE10", X"0270", X"0046", X"FF00", X"FEFC", X"FED8", X"FF06", X"011F", X"0449", X"073D", X"0755", X"0787", X"06F9", X"0072", X"01C0", X"015D", X"0149", X"0011", X"FF7A", X"FF3F", X"00A3", X"FF42", X"FF5E", X"006A", X"01E3", X"FBF5", X"F963", X"FD44", X"FE0B", X"FF04", X"00B0", X"03D7", X"0129", X"FFB3", X"0133", X"026D", X"0344", X"0507", X"0580", X"0518", X"03E8", X"00C3", X"01A0", X"0249", X"00AA", X"0249", X"0473", X"0171", X"0019", X"FD8C", X"FE9B", X"FD22", X"FB9A", X"F8D2", X"FBD2", X"FD29", X"FB36", X"FF0E", X"027C", X"0223", X"FF90", X"FED1", X"0038", X"FE99", X"FEDB", X"00D4", X"0481", X"03A9", X"02EA", X"06F0", X"04DD", X"0614", X"04C3", X"0645", X"03BA", X"01A0", X"FFBF", X"005E", X"FF5B", X"0152", X"FF3D", X"FC76", X"FB48", X"FB72", X"FCEB", X"0198", X"FE39", X"0050", X"FECC", X"FFE4", X"FF92", X"0071", X"FDF4", X"FD7C", X"0033", X"010E", X"0108", X"03D4", X"0164", X"006A", X"0119", X"0154", X"FFDE", X"00EA", X"023B", X"03DD", X"04A0", X"0554", X"067A", X"003C", X"FDFB", X"FF17", X"FDE1", X"0043", X"00A1", X"FF8D", X"010F", X"FEC1", X"007D", X"00F3", X"FEC2", X"006E", X"02F6", X"00AC", X"01E9", X"024D", X"02AE", X"025B", X"004D", X"0147", X"07FA", X"044A", X"0266", X"05C5", X"066B", X"0457", X"051F", X"012A", X"FFA0", X"FF88", X"0161", X"FF6C", X"FFAF", X"01BA", X"FF5A"),
        (X"00DC", X"01A6", X"00E3", X"FF1F", X"FF17", X"0124", X"000E", X"FF8A", X"FDE9", X"0100", X"015B", X"FFBE", X"00F1", X"00CB", X"00CA", X"FEAA", X"00D6", X"FFEE", X"FEC0", X"FFCF", X"FF89", X"01DB", X"00DB", X"0055", X"00FF", X"004B", X"FF0F", X"0055", X"FF43", X"00FC", X"0078", X"00E3", X"0059", X"00ED", X"0374", X"03C6", X"01C6", X"025A", X"03E7", X"0592", X"03E0", X"02CB", X"FF8F", X"0498", X"02CF", X"00DA", X"0445", X"0401", X"03C7", X"02BF", X"02CA", X"022B", X"FFDB", X"008C", X"FFEA", X"FFFB", X"FDE5", X"014A", X"0131", X"00C0", X"01BB", X"00C8", X"0308", X"04A0", X"06C0", X"0956", X"078D", X"0B01", X"0A95", X"04DF", X"0692", X"0519", X"0558", X"03B2", X"0612", X"061E", X"0682", X"05CA", X"039C", X"04F8", X"0342", X"0107", X"00D8", X"FF20", X"01FE", X"FFE8", X"00BC", X"0162", X"0172", X"0750", X"05C8", X"05EF", X"0807", X"09B8", X"078B", X"0674", X"0973", X"08EA", X"05C4", X"030A", X"00D2", X"0213", X"035A", X"0077", X"0339", X"041B", X"0330", X"0737", X"05E0", X"0390", X"0115", X"0069", X"00FB", X"FFF3", X"FFD1", X"00D4", X"0279", X"0509", X"051E", X"0359", X"045F", X"04CF", X"06E8", X"041C", X"0442", X"039F", X"041F", X"0372", X"0309", X"02FB", X"044E", X"03C3", X"03AE", X"034E", X"0259", X"0135", X"01E6", X"FF7D", X"0208", X"0165", X"FFB5", X"FF7F", X"016C", X"01B4", X"051C", X"02E8", X"0271", X"03E9", X"0357", X"0170", X"013F", X"FF8A", X"FE51", X"FE3D", X"FF88", X"020C", X"02A7", X"037A", X"0403", X"02D6", X"0253", X"0076", X"FF9C", X"01CD", X"01F3", X"00C7", X"00DB", X"031D", X"FE4F", X"0112", X"FD66", X"02DB", X"022E", X"017F", X"006E", X"01FE", X"017D", X"0279", X"000E", X"FFDE", X"005E", X"0192", X"019B", X"031F", X"026F", X"0050", X"0025", X"FE56", X"FF08", X"FE24", X"FD3D", X"FE66", X"FED8", X"FFFE", X"FEF6", X"017E", X"FFE8", X"0240", X"002F", X"FFFA", X"03E2", X"0174", X"00DF", X"FE98", X"0025", X"FF57", X"0094", X"FFE7", X"0356", X"01E1", X"0247", X"01BD", X"FFAD", X"FCFB", X"FCBA", X"FD24", X"FCBD", X"FCC9", X"FC18", X"F816", X"FB0A", X"FCA4", X"FFF0", X"027D", X"FE24", X"0105", X"FCB8", X"FF63", X"03DC", X"FF5B", X"FDD8", X"FD59", X"FE68", X"FEFA", X"00E6", X"FFE1", X"0267", X"039F", X"0201", X"FD2D", X"FC8A", X"F9C3", X"F875", X"FBF9", X"FC2C", X"FD22", X"FCA1", X"F7AB", X"F431", X"F768", X"FB1A", X"FCB9", X"003E", X"FDC4", X"0150", X"0062", X"041A", X"FC72", X"FBAF", X"FE38", X"FFD0", X"FDF0", X"FD47", X"FECE", X"0059", X"0031", X"00A9", X"FE8D", X"FAE2", X"F852", X"F9AC", X"FB63", X"FDB7", X"FDA5", X"FE6D", X"FB7C", X"F6F9", X"F82E", X"FD1A", X"0098", X"001A", X"FF51", X"00B5", X"0299", X"FF91", X"FD0F", X"FD6B", X"FD19", X"FC66", X"FA44", X"FA31", X"FC34", X"FC80", X"FF81", X"032B", X"01DE", X"FCD7", X"FACF", X"F9E2", X"FCDC", X"003B", X"FEB9", X"FD5C", X"FE1C", X"FB9E", X"FBED", X"FCF4", X"FCA2", X"008D", X"FE35", X"0090", X"0395", X"FF2E", X"FC7F", X"F94F", X"F87B", X"F8C6", X"F983", X"F86F", X"FB2E", X"FAA8", X"0071", X"048C", X"0311", X"FFCD", X"FC6C", X"FE02", X"0001", X"FE9D", X"FC37", X"FE8C", X"005F", X"014F", X"0052", X"FBBB", X"FEC5", X"FFE6", X"FD8C", X"FD62", X"FDBE", X"FCE2", X"FA37", X"F7D2", X"F7B2", X"FBE0", X"FAB4", X"FB46", X"F9F8", X"FB45", X"010A", X"0700", X"03F9", X"02E2", X"FF21", X"FF36", X"FCD9", X"FDF5", X"FE89", X"FE0E", X"FEE7", X"0244", X"0269", X"FDD9", X"0280", X"FF75", X"FDE8", X"FD70", X"008E", X"FBFE", X"F9C4", X"FB68", X"F99F", X"FBBF", X"FC2A", X"FB94", X"FA2D", X"FC3B", X"0432", X"05B7", X"0415", X"0183", X"026E", X"FEA8", X"FCEB", X"FB06", X"FD95", X"FD9F", X"0177", X"02F4", X"0265", X"027B", X"02F6", X"FEDB", X"FF38", X"FC84", X"016B", X"FAB3", X"FD88", X"004E", X"FCEA", X"FD47", X"FD32", X"FA21", X"FD23", X"FD35", X"031F", X"07AD", X"06A9", X"0298", X"FF0E", X"0004", X"FE79", X"FF29", X"0066", X"0054", X"00E3", X"0284", X"025A", X"07B7", X"03BB", X"FDCB", X"00EA", X"022A", X"02B9", X"FE0B", X"0024", X"00EA", X"FF92", X"FDCD", X"FD6B", X"FC9F", X"FFA7", X"0220", X"0612", X"06E3", X"05CE", X"0212", X"FF28", X"FF79", X"FEC4", X"0015", X"0074", X"002B", X"0078", X"031E", X"058F", X"059C", X"018A", X"FFD3", X"0054", X"048B", X"068C", X"00FE", X"FF24", X"FEE0", X"FD33", X"FB82", X"FE49", X"00DC", X"029B", X"061C", X"05EC", X"0312", X"037A", X"FF59", X"00F0", X"0295", X"0317", X"02C3", X"0146", X"01FD", X"0134", X"056D", X"084D", X"0660", X"0344", X"FFF0", X"01C1", X"03A0", X"06A6", X"00DD", X"FFEC", X"0006", X"00DC", X"FD2E", X"FE21", X"FE9C", X"02BF", X"01D1", X"01B1", X"01C6", X"0108", X"0070", X"00DB", X"036A", X"040D", X"0367", X"01B5", X"02FB", X"01E8", X"0117", X"077C", X"04AF", X"FFB8", X"FFAF", X"0183", X"0024", X"0771", X"020E", X"01D4", X"0083", X"002E", X"FF4E", X"FF51", X"0042", X"025D", X"000C", X"011E", X"FED8", X"010C", X"0353", X"03A6", X"0420", X"01E7", X"01A3", X"02DA", X"028C", X"034D", X"0176", X"0876", X"0452", X"0322", X"00FB", X"FD2E", X"FF11", X"0604", X"02FB", X"01E8", X"00E1", X"00CE", X"0103", X"0373", X"03C1", X"04CE", X"00A0", X"0044", X"0051", X"02A4", X"0623", X"04CB", X"01AC", X"030C", X"02E6", X"0350", X"0249", X"0077", X"0265", X"0564", X"03F5", X"015C", X"00D2", X"FBEA", X"001A", X"0760", X"065D", X"02CD", X"02E8", X"0316", X"0407", X"048B", X"0445", X"00E9", X"FF41", X"FEF9", X"00BB", X"03BE", X"043C", X"02B0", X"0167", X"01A5", X"03C0", X"017B", X"0061", X"FFAC", X"0283", X"0129", X"029A", X"FF74", X"FFD2", X"008A", X"0417", X"0804", X"033D", X"01F1", X"0109", X"0284", X"051E", X"040C", X"02CB", X"0218", X"FE7B", X"00B9", X"0344", X"024B", X"0518", X"021C", X"01FA", X"01BF", X"01A5", X"FF15", X"FF96", X"00AF", X"00A6", X"0064", X"FF50", X"FF30", X"FFEC", X"FEB4", X"0374", X"0818", X"0513", X"0241", X"0079", X"0120", X"0087", X"010E", X"0142", X"FE82", X"FE2E", X"FEE1", X"FEBC", X"0104", X"0145", X"00E8", X"FF75", X"0241", X"017A", X"00CA", X"FDA1", X"FF7B", X"FBEF", X"FF49", X"FE3B", X"0005", X"0187", X"00C2", X"047E", X"06C0", X"05FD", X"03B6", X"02CE", X"0267", X"0205", X"FF6D", X"FEA2", X"FE2E", X"FB90", X"FCD6", X"FD60", X"FFDE", X"FEBB", X"01A5", X"007F", X"0114", X"00B8", X"FF05", X"FFE2", X"FEAA", X"FBE8", X"FE08", X"0185", X"FF7B", X"FFD6", X"009C", X"00A0", X"018E", X"031C", X"007A", X"0271", X"0453", X"02D7", X"01A1", X"00EF", X"FF01", X"FF2A", X"FEAD", X"FEC3", X"FED0", X"FFFF", X"019D", X"01ED", X"FE15", X"FF27", X"FE56", X"FF7A", X"FEB6", X"03F6", X"0454", X"0202", X"00AE", X"00C8", X"0088", X"0125", X"FC37", X"FD6A", X"0072", X"0243", X"0376", X"0683", X"052F", X"0258", X"03D2", X"048A", X"029C", X"0197", X"FE81", X"03A6", X"04E9", X"044D", X"032A", X"006D", X"FF51", X"FE67", X"FD19", X"0016", X"0249", X"01A8", X"FF31", X"FF52", X"00A4", X"FF4D", X"FFEB", X"FCC7", X"FFCA", X"FE98", X"FF06", X"FDB2", X"FE71", X"FC1D", X"FD8C", X"0158", X"FFE6", X"0081", X"FFDE", X"04B8", X"0373", X"0486", X"0227", X"03A9", X"FFB9", X"FE5F", X"0046", X"FFDF", X"FFD0", X"012D", X"FF57", X"00AF", X"FFA1", X"FFCC", X"0006", X"016C", X"0107", X"00B2", X"FF1A", X"00C2", X"FED2", X"003A", X"01F3", X"FF68", X"FF08", X"FE4B", X"FB90", X"FB5E", X"FC1E", X"FCF9", X"FD01", X"FF2D", X"FE9B", X"FDF6", X"FFE8", X"00E2", X"FF79", X"0047", X"FF3F"),
        (X"006E", X"FEA8", X"012A", X"FF39", X"FFD2", X"FEA8", X"0006", X"001A", X"0029", X"FF08", X"FFC0", X"0052", X"0092", X"0138", X"0053", X"FFDF", X"0020", X"0158", X"00CE", X"FFDD", X"00F1", X"0030", X"00BB", X"FEEF", X"FFBA", X"00B5", X"0013", X"014E", X"FEFE", X"FFE8", X"006B", X"FF83", X"0042", X"0017", X"005A", X"FF38", X"FF66", X"FF76", X"FE0C", X"01CD", X"01EC", X"01F6", X"FCAC", X"0176", X"01BE", X"012C", X"FD77", X"FBEB", X"FF17", X"FF8A", X"0078", X"027F", X"FF20", X"0022", X"FF47", X"FF57", X"FFD6", X"FF62", X"0024", X"01AD", X"0188", X"FF8C", X"FE75", X"FFB5", X"FE13", X"FD91", X"FD01", X"FBF5", X"FE3F", X"FADC", X"F4AB", X"F574", X"F9EC", X"F9EC", X"FD48", X"FC97", X"FBDF", X"F8F2", X"F9AA", X"FB00", X"00F9", X"015F", X"006F", X"FF8B", X"FEDF", X"FF05", X"0017", X"0061", X"00BB", X"FB6D", X"FBA8", X"FAED", X"FB38", X"FC86", X"FBC1", X"F9E6", X"F9A1", X"FA24", X"FAF8", X"F8AD", X"F862", X"F890", X"F91C", X"FAE1", X"FC31", X"FED9", X"FE92", X"FE33", X"FFB9", X"01BD", X"FEB5", X"FEEF", X"00CF", X"004F", X"FDD6", X"0147", X"FAF4", X"F721", X"FAE3", X"FC11", X"F89E", X"FC43", X"FBB9", X"FCE9", X"FA2B", X"F941", X"FB48", X"FC6F", X"FA57", X"FBFA", X"FB18", X"FC1D", X"FCFE", X"FF80", X"FF7D", X"012B", X"00E4", X"02DE", X"0382", X"FD89", X"FF23", X"FFEF", X"FDA9", X"FDFA", X"F91A", X"F8AF", X"FC7D", X"FD06", X"FDFC", X"FC50", X"FE17", X"0019", X"FE3E", X"00C0", X"002B", X"FD57", X"FDDF", X"00B7", X"00F6", X"FFAD", X"015E", X"0103", X"00BA", X"FD24", X"FEB8", X"0168", X"FFD3", X"FE9B", X"0074", X"FF54", X"FE5B", X"FD8F", X"FAE8", X"FD96", X"FECA", X"FE4E", X"FD7B", X"FC77", X"FE81", X"FE71", X"024A", X"03F8", X"03F8", X"050A", X"050C", X"05CA", X"059F", X"0309", X"0108", X"00B8", X"FF70", X"00D8", X"02D7", X"0225", X"00AC", X"FFC4", X"00B8", X"FEE3", X"007B", X"FDAC", X"F999", X"FB96", X"FDCC", X"FC28", X"FE4D", X"FDAC", X"0196", X"0403", X"04BF", X"05B9", X"04F6", X"050B", X"063E", X"03CB", X"02AC", X"0094", X"FF55", X"00D2", X"00AC", X"069A", X"0AA6", X"0A46", X"0419", X"FF8C", X"0283", X"01F3", X"011E", X"FFC9", X"FB6E", X"FCA5", X"FDF2", X"FEA1", X"0320", X"0338", X"04C6", X"05C2", X"0598", X"048A", X"054E", X"036C", X"02AF", X"01A9", X"000B", X"00F4", X"FF82", X"01CE", X"04E7", X"0C2E", X"1071", X"0EE3", X"05A7", X"0367", X"017C", X"01AF", X"0244", X"0135", X"FCC5", X"FE7B", X"01D0", X"039F", X"05AB", X"0605", X"0895", X"080F", X"062C", X"05BF", X"0493", X"00BF", X"0009", X"00CD", X"0134", X"004C", X"0063", X"033C", X"079A", X"0DEB", X"12D6", X"0D29", X"088A", X"03FB", X"FE86", X"0224", X"0482", X"01E6", X"019A", X"03D4", X"057D", X"04F9", X"07F8", X"072D", X"0720", X"04F0", X"0467", X"03ED", X"02A4", X"FF27", X"FED7", X"0024", X"00C9", X"0109", X"0296", X"06FA", X"0B35", X"0DDE", X"0D6D", X"0C55", X"0673", X"022B", X"00CD", X"02FE", X"05E7", X"0319", X"0577", X"0896", X"0907", X"0942", X"08BC", X"0409", X"00B7", X"0275", X"00D4", X"03F5", X"FE94", X"FD8E", X"FE42", X"00F7", X"019F", X"00DF", X"06CC", X"078C", X"09E5", X"09C2", X"08E3", X"08E1", X"05A1", X"01D7", X"001F", X"00BD", X"0658", X"05BC", X"0849", X"09A3", X"066C", X"03FD", X"0169", X"FEE6", X"FE3A", X"FC97", X"FA85", X"FB1D", X"FBC4", X"FD58", X"FDBF", X"009B", X"016B", X"02E5", X"0302", X"03A7", X"027A", X"FE01", X"FA90", X"FF66", X"0288", X"030C", X"FFAF", X"0179", X"044D", X"05C5", X"05A0", X"0305", X"02CE", X"0126", X"FCD5", X"FD88", X"FD24", X"FB5C", X"FC3C", X"FCB2", X"FCD0", X"FB65", X"FD15", X"FF78", X"0099", X"FFAD", X"0195", X"FF64", X"00DD", X"FBEB", X"FA5B", X"FDCE", X"FF33", X"00AC", X"0113", X"01C2", X"03FD", X"0180", X"FD03", X"FD1F", X"FD5D", X"FE6A", X"FD0A", X"FD24", X"FF3C", X"FEF0", X"FBDC", X"FCB2", X"F9D6", X"FD3B", X"FC83", X"FEBE", X"FE8B", X"FE0F", X"FFAB", X"FDB2", X"FCE4", X"FB95", X"FD2F", X"FCDD", X"019C", X"027F", X"0234", X"FDAF", X"FC46", X"FA34", X"FC02", X"FB47", X"FC9C", X"FC70", X"FC35", X"FED4", X"FF27", X"FFDB", X"FD3B", X"FBB9", X"F7A3", X"FAC3", X"FD0B", X"004B", X"0110", X"FEFE", X"FF89", X"FF32", X"FC98", X"FC7B", X"FFCC", X"FBFD", X"FC59", X"FEF8", X"01F5", X"FCB4", X"FAA4", X"F87A", X"FDAA", X"FDA1", X"FC57", X"FA90", X"FA24", X"FD47", X"0054", X"0006", X"FE28", X"FB3C", X"FA06", X"FD1C", X"FDDC", X"0088", X"FF29", X"FCFF", X"FD13", X"FC49", X"FDA6", X"FB06", X"FA87", X"FA2F", X"FDA4", X"FDB1", X"FFB2", X"FD86", X"F92A", X"F8B4", X"FD08", X"0248", X"01C5", X"FC9E", X"FDCE", X"FF03", X"FFCE", X"0178", X"FEA4", X"FC36", X"FCC1", X"FEF2", X"00CA", X"FE9B", X"FDAF", X"FE40", X"FD28", X"FAC2", X"FBE7", X"FC00", X"FD43", X"FEC3", X"FEBD", X"FFFE", X"0313", X"005A", X"FBFE", X"F6B0", X"FE48", X"0186", X"01DC", X"0300", X"0135", X"0081", X"01D8", X"02BC", X"FE9B", X"FFF2", X"0044", X"0040", X"FEBC", X"000E", X"FDEE", X"FE5B", X"FB7D", X"FBCB", X"FCEB", X"FC40", X"FEFC", X"0050", X"FD5D", X"FC02", X"FF71", X"0376", X"00E5", X"F4CB", X"FF41", X"0122", X"021C", X"0126", X"0203", X"01F8", X"03A9", X"0297", X"03ED", X"0179", X"0172", X"FD99", X"FD4A", X"FCBA", X"FBF7", X"FEA6", X"FC5A", X"FC4A", X"FEEB", X"030A", X"0676", X"0457", X"FD1C", X"FEAD", X"00CB", X"02BF", X"FE96", X"F9F4", X"FF51", X"03F7", X"0165", X"013A", X"00AC", X"01DA", X"0251", X"018C", X"00F6", X"FFE9", X"FE86", X"FD45", X"FD37", X"FF2C", X"FD40", X"FE8C", X"FC1D", X"FD62", X"01F8", X"05D2", X"0984", X"063C", X"FD15", X"FF2B", X"FFC5", X"FD83", X"FC72", X"FAA9", X"0061", X"0208", X"0448", X"040A", X"022F", X"02BB", X"0115", X"FF5E", X"FF64", X"FF8D", X"FCCD", X"FC1F", X"FD8F", X"FCB9", X"FC96", X"FC71", X"FC0E", X"FF55", X"03D1", X"0563", X"072D", X"0574", X"0151", X"FFEF", X"0180", X"FF99", X"FC2E", X"FAD6", X"01D2", X"00F3", X"03CC", X"065B", X"054A", X"0340", X"0136", X"00DC", X"019B", X"0002", X"0146", X"FF89", X"FFC7", X"FF3C", X"FE6B", X"FD2A", X"FC61", X"FF8F", X"03F6", X"07EC", X"0703", X"0535", X"0291", X"FE9B", X"FF9F", X"00CE", X"FBD5", X"FB6E", X"FE8E", X"FF36", X"0036", X"0185", X"02AC", X"0264", X"0300", X"01AF", X"01F3", X"012E", X"FFD2", X"FFB9", X"019E", X"016E", X"FDEA", X"FFB3", X"0103", X"0133", X"0243", X"0611", X"05E7", X"0318", X"FD20", X"001E", X"00B6", X"0019", X"0155", X"FC0D", X"FE98", X"FFFE", X"FF77", X"FE52", X"FF9D", X"FE2C", X"FF56", X"FDD3", X"008B", X"FF41", X"007C", X"02CC", X"02CB", X"035A", X"0369", X"0417", X"0390", X"02B0", X"017A", X"04C3", X"02AE", X"FD62", X"FD63", X"002A", X"0050", X"FF8E", X"0020", X"FFE2", X"015A", X"0188", X"01D1", X"0239", X"0187", X"01AA", X"00CF", X"0315", X"027F", X"01C9", X"0421", X"0570", X"0683", X"06E1", X"0795", X"06FA", X"076B", X"050C", X"0469", X"0225", X"037A", X"FE96", X"FEB4", X"FE77", X"FE5D", X"FF86", X"0046", X"00C4", X"03D4", X"0757", X"08A8", X"063C", X"0B51", X"0E4C", X"0D2E", X"0CDA", X"0D27", X"0F75", X"1127", X"0BC5", X"0B02", X"0AA0", X"0B08", X"0738", X"08E6", X"0768", X"0503", X"02DC", X"015C", X"FFAC", X"FEDA", X"00C2", X"0094", X"00E3", X"FF02", X"FEC3", X"00BA", X"01D3", X"0454", X"0452", X"03C4", X"05D2", X"0810", X"04A8", X"0752", X"0756", X"095A", X"0562", X"04EB", X"06EF", X"0662", X"026F", X"025D", X"02C7", X"00E6", X"01CA", X"FF9F", X"FEA7", X"0051", X"0084"),
        (X"0049", X"FEE4", X"FFE1", X"0137", X"FE69", X"FFB3", X"FFB6", X"00A4", X"0009", X"012F", X"0020", X"00E7", X"008E", X"FF3B", X"FFF6", X"FFEC", X"FFD8", X"00EE", X"016C", X"FED0", X"00E0", X"0037", X"FF90", X"0075", X"FDE1", X"0099", X"0234", X"0051", X"FFDA", X"00D8", X"020B", X"FF12", X"008A", X"FEEC", X"FE8D", X"FE52", X"FFC2", X"FEFC", X"FF50", X"01BA", X"027B", X"0085", X"FD0B", X"FECA", X"003F", X"00C4", X"FD9B", X"FE97", X"FF1C", X"FEE0", X"0030", X"FFDB", X"00F2", X"FFF6", X"FFBD", X"FFC1", X"FE52", X"00AE", X"003A", X"0202", X"0281", X"0002", X"FD3A", X"FF70", X"FC9B", X"F764", X"F8A1", X"FA8F", X"FBCD", X"FB56", X"F839", X"F921", X"FFEA", X"0089", X"FEF2", X"015F", X"FED9", X"FD4F", X"FFAF", X"FE01", X"FDDC", X"0075", X"FF12", X"FFCA", X"00AE", X"FFB3", X"00DA", X"00FF", X"019B", X"024C", X"FF7A", X"FE75", X"0052", X"FCDA", X"FF20", X"012A", X"012D", X"FFF7", X"0220", X"02D5", X"048D", X"0492", X"00E8", X"0134", X"0196", X"008D", X"FCB4", X"FB09", X"FC0E", X"FF82", X"0164", X"FFE9", X"00C8", X"FFED", X"02A9", X"0423", X"FF42", X"FE93", X"FD16", X"FD1B", X"FC54", X"FBF0", X"FCCA", X"FF89", X"FDF8", X"FC09", X"FF42", X"FEE2", X"FFE5", X"FF18", X"FFFA", X"FE6D", X"FC6F", X"FD60", X"FE68", X"FE16", X"FFD0", X"01B8", X"00A7", X"FD75", X"FF55", X"00E5", X"FD32", X"0076", X"FE14", X"007F", X"FF4B", X"0097", X"01FC", X"FF49", X"0067", X"000C", X"00BF", X"00FE", X"0151", X"0073", X"FF4D", X"FE22", X"FE40", X"FF0B", X"FD8A", X"FCCE", X"FFB9", X"FED4", X"FE80", X"02BB", X"025C", X"FCCD", X"0061", X"0091", X"01A0", X"0331", X"01E0", X"0643", X"04A8", X"0668", X"0502", X"05DC", X"0783", X"050D", X"0456", X"056A", X"02CB", X"0115", X"0092", X"FF67", X"0111", X"FFC9", X"00A4", X"007E", X"015E", X"FF1C", X"0263", X"FF78", X"FF72", X"01D2", X"003D", X"0438", X"FFE4", X"05A6", X"0522", X"0832", X"066B", X"0728", X"0509", X"0691", X"05A8", X"05FE", X"046C", X"041B", X"FFD3", X"0136", X"0269", X"0325", X"00FE", X"0076", X"0386", X"0183", X"0203", X"027E", X"0122", X"03EE", X"0167", X"0119", X"01AE", X"02AB", X"0104", X"05E8", X"04A4", X"0627", X"06E7", X"04D7", X"0360", X"030A", X"058B", X"0485", X"03BD", X"026B", X"021D", X"0244", X"014B", X"0382", X"0428", X"02F5", X"026F", X"0119", X"02D8", X"04C6", X"0580", X"0436", X"0275", X"01D3", X"00B8", X"0419", X"03A3", X"06B4", X"055C", X"04B4", X"01E7", X"015D", X"00B1", X"01C7", X"00B1", X"0333", X"017F", X"005C", X"03F1", X"0439", X"0425", X"045B", X"03CE", X"03F0", X"0256", X"01C6", X"032B", X"043A", X"07D7", X"07D1", X"0527", X"026B", X"01E1", X"0355", X"05D6", X"0713", X"030C", X"03D1", X"FE17", X"FDAF", X"FE63", X"FF2A", X"FFAA", X"0147", X"02D6", X"02DC", X"0462", X"059B", X"06D8", X"046A", X"0355", X"011D", X"0322", X"00E3", X"0167", X"0380", X"06F3", X"09D1", X"09D9", X"01DB", X"FFCD", X"0480", X"0637", X"05E7", X"019C", X"FD23", X"FEB3", X"FD62", X"FC86", X"FC73", X"FE55", X"0302", X"0514", X"05FC", X"0566", X"0690", X"0492", X"0422", X"008B", X"FD62", X"FD9F", X"FB7A", X"FCBD", X"FE4E", X"FF47", X"063E", X"04E3", X"0141", X"01E5", X"0581", X"070D", X"038F", X"FD41", X"FDA5", X"FC5B", X"FC84", X"FE44", X"FB40", X"FCE7", X"001B", X"009A", X"01EC", X"0063", X"000F", X"FEA9", X"FE5F", X"FD69", X"FA3D", X"F999", X"F815", X"F8C9", X"FBD1", X"FEF0", X"FF9D", X"0222", X"FDEA", X"FFFE", X"02F3", X"06E3", X"FFBC", X"FC69", X"FB59", X"FDCE", X"FB46", X"FA73", X"FC2C", X"FA27", X"F902", X"F8E4", X"F863", X"FB1F", X"FAB6", X"FDAB", X"FF55", X"FDB2", X"FAA3", X"FB7A", X"FAA4", X"FC79", X"FFB1", X"02A1", X"FEBF", X"FBEC", X"FF06", X"0286", X"0330", X"0637", X"0078", X"FC8F", X"FE42", X"FBB1", X"FD14", X"FB47", X"FB11", X"FAFD", X"F589", X"F63D", X"F54C", X"F8DE", X"FA22", X"FBEC", X"002C", X"01AA", X"01E9", X"010B", X"FF7D", X"038F", X"0777", X"0788", X"FCA1", X"FB2E", X"FCC8", X"015F", X"02A3", X"03C1", X"FEDE", X"FE1D", X"FEA1", X"FD80", X"FB89", X"FD43", X"FD2B", X"FD4B", X"FBE8", X"FC19", X"F973", X"F7F4", X"FC12", X"FB52", X"0094", X"02A3", X"0496", X"0503", X"0730", X"05E0", X"06D7", X"06A1", X"F988", X"F931", X"FCF2", X"01CA", X"0124", X"0369", X"0012", X"016C", X"FE16", X"FD6F", X"FC60", X"FEFA", X"FE19", X"FE29", X"FD92", X"FD8F", X"FC7D", X"FB2B", X"FB53", X"FC66", X"FF1D", X"01B7", X"044B", X"059A", X"03AC", X"03E8", X"04A8", X"0381", X"F54A", X"F725", X"FE09", X"FF77", X"0201", X"017F", X"01E8", X"0382", X"FFDE", X"FE6A", X"FC40", X"FC0A", X"FC8B", X"FC7B", X"FC51", X"FB83", X"FBF3", X"FBA4", X"FBFB", X"FD73", X"029D", X"0468", X"0353", X"0391", X"0457", X"0247", X"026F", X"0207", X"FB7F", X"FF6D", X"0169", X"0136", X"0131", X"0394", X"04B6", X"02BC", X"02CC", X"FEBA", X"F975", X"FC97", X"F9B5", X"FA22", X"FBE4", X"FAC4", X"FAAC", X"FCBD", X"FE86", X"FEAE", X"0223", X"0307", X"0258", X"011C", X"0178", X"021A", X"FF2D", X"FD8A", X"FA41", X"0039", X"FB9E", X"00D5", X"0396", X"03EE", X"05AD", X"0571", X"0354", X"FFFE", X"FBCF", X"FEF4", X"FE7C", X"FCEB", X"FE59", X"FF7A", X"FD7A", X"FE86", X"FD63", X"FD2A", X"00F2", X"FF81", X"FED6", X"FDE3", X"FDD7", X"FDF8", X"FBD3", X"FC77", X"F851", X"FB89", X"FF33", X"FFBF", X"037A", X"0264", X"0542", X"0108", X"0196", X"FF8F", X"FD57", X"004D", X"0153", X"03BA", X"034F", X"02C6", X"00B8", X"007E", X"FDE6", X"FE22", X"FE96", X"FE52", X"FC5F", X"FA52", X"FC51", X"FDB4", X"FAE8", X"F916", X"FA13", X"FECD", X"004D", X"00B1", X"FEA8", X"025B", X"036A", X"0045", X"FFCC", X"01A2", X"FFF9", X"FFA9", X"0196", X"023F", X"0266", X"0345", X"00B7", X"0005", X"00F5", X"00CC", X"FF4B", X"FE44", X"FC20", X"FA77", X"FBF2", X"FC85", X"F818", X"F600", X"F911", X"FFB3", X"FF17", X"FE91", X"FE7F", X"030D", X"0353", X"FFE8", X"0164", X"00A6", X"009A", X"0233", X"002F", X"0190", X"026E", X"02F4", X"01DC", X"01BF", X"0241", X"017E", X"01CE", X"FF33", X"FD7E", X"FAF1", X"FC07", X"FBE4", X"F723", X"F5F3", X"FA6A", X"FEC1", X"0161", X"FFC4", X"FFB5", X"0332", X"04B8", X"0662", X"0662", X"05D4", X"0796", X"025B", X"02A4", X"02B0", X"03F0", X"0369", X"0401", X"028C", X"0359", X"036B", X"0104", X"FD3A", X"F995", X"F73E", X"F72E", X"F97D", X"F55E", X"F727", X"FC0B", X"FFCC", X"003A", X"FF65", X"FF53", X"008C", X"04EE", X"0A65", X"0B27", X"08D8", X"06AB", X"034F", X"0571", X"04B6", X"023F", X"04E0", X"05A3", X"0495", X"03C1", X"0069", X"FF6E", X"FC0E", X"FA3F", X"F7DB", X"F81F", X"F958", X"FA1F", X"FC39", X"FB57", X"FFDE", X"FF14", X"FFDF", X"FFD4", X"FE78", X"033E", X"05EF", X"0570", X"0350", X"0260", X"0390", X"0584", X"0338", X"0447", X"03B1", X"02EC", X"FF56", X"FFF7", X"FE7B", X"FFA6", X"0130", X"0162", X"FA41", X"FBF7", X"FF9A", X"FCE5", X"0099", X"FFB8", X"FF60", X"006B", X"FF84", X"FE6D", X"000F", X"FF76", X"FC32", X"FF07", X"FCAB", X"FBFA", X"FE7B", X"FFAD", X"0024", X"FDDD", X"FC81", X"FF08", X"FD8E", X"0081", X"0048", X"01C1", X"031E", X"049A", X"013E", X"FDC5", X"003E", X"FEB4", X"FE95", X"0131", X"0090", X"FFBD", X"FFC4", X"0050", X"0053", X"0026", X"0155", X"015B", X"0091", X"FE22", X"009D", X"0193", X"0368", X"0168", X"01DF", X"061D", X"0174", X"00D8", X"01B9", X"0537", X"0116", X"051B", X"0130", X"018A", X"00A9", X"03FA", X"FFDB", X"00F7", X"0135", X"FFE6"),
        (X"0063", X"FF89", X"FF79", X"FF04", X"FF6D", X"FE7A", X"001A", X"FEC1", X"001B", X"FEBD", X"00E9", X"FF35", X"FF58", X"FDF4", X"0016", X"FF9B", X"005A", X"0044", X"FF3F", X"FFFD", X"FEC5", X"0099", X"FFB0", X"0129", X"00C7", X"FEE2", X"FEFD", X"008B", X"0168", X"FF5C", X"0000", X"FE99", X"FEA6", X"FF96", X"FAF6", X"FC1F", X"FC26", X"FA47", X"F9F5", X"FA86", X"F9C1", X"FC24", X"00DF", X"00C0", X"FC3C", X"FA97", X"FC2B", X"FCF3", X"F8B3", X"FDE7", X"FE00", X"FD51", X"FF3D", X"006C", X"FF56", X"FFD7", X"FF69", X"FFDB", X"0001", X"FCD5", X"FCCF", X"FE11", X"F9EF", X"F9F0", X"F75A", X"F4F2", X"F59E", X"F48C", X"F610", X"F92B", X"FCB7", X"FCC3", X"FC5D", X"FD77", X"F9C9", X"F735", X"F90F", X"F9A3", X"F9E1", X"F885", X"FBA9", X"FDC6", X"00F4", X"FF20", X"FF09", X"00AD", X"027D", X"FC71", X"FDE1", X"010B", X"FAAB", X"F78C", X"F889", X"F8FB", X"FC25", X"FE89", X"FFB3", X"FE69", X"000C", X"FF9A", X"0016", X"FF3F", X"FDD7", X"FCF2", X"FFEC", X"F982", X"F86E", X"F79E", X"F8CF", X"FB8D", X"FD3C", X"0103", X"FF77", X"FF82", X"00CE", X"03D5", X"05DB", X"06E9", X"04CC", X"03FB", X"026B", X"FE0D", X"FE4D", X"0021", X"FF60", X"00BC", X"FF77", X"FEBB", X"FDAB", X"FD7E", X"FE81", X"FF13", X"FE95", X"FF14", X"005C", X"FDCF", X"FAC3", X"F9EA", X"FC03", X"FCD8", X"0064", X"FFDC", X"017C", X"048B", X"0726", X"0A93", X"07BF", X"0396", X"FEDD", X"FF50", X"FD57", X"FDC5", X"FE8A", X"FC6A", X"FCEA", X"FF89", X"FD7A", X"FD28", X"FCF9", X"FD18", X"FCD5", X"FDB0", X"FE1E", X"FE47", X"FA3B", X"F4CA", X"FA2D", X"FEE2", X"FFE5", X"FF31", X"0045", X"075C", X"09E6", X"0925", X"0602", X"02F7", X"00C7", X"01B6", X"FFD0", X"FEDD", X"FEE9", X"FE02", X"FF0F", X"FDE2", X"007F", X"00FB", X"0273", X"006E", X"FF06", X"FF07", X"FF85", X"FE13", X"F8A6", X"F4FD", X"FB9B", X"FD81", X"0023", X"01F8", X"FFD0", X"0786", X"0B88", X"0803", X"03B8", X"01A9", X"FDF2", X"FE87", X"FE2A", X"FF52", X"FF41", X"FF44", X"00B5", X"021F", X"0377", X"049E", X"01B9", X"02A9", X"01F4", X"FF25", X"0018", X"FBE3", X"F628", X"F37B", X"FAAC", X"FC36", X"FEB6", X"FEEB", X"00F8", X"0485", X"07F7", X"02FA", X"0173", X"008A", X"FFAA", X"FE78", X"FD04", X"FD3D", X"FBF8", X"FEC7", X"037D", X"0599", X"0555", X"0503", X"0549", X"03BC", X"03DD", X"03F7", X"FFC0", X"FB1F", X"F5A0", X"F846", X"F855", X"FEDE", X"0049", X"02D1", X"00BD", X"0135", X"052A", X"013F", X"02C8", X"005A", X"FE14", X"FCA5", X"FAA6", X"F970", X"FA09", X"FDC6", X"04F9", X"08EB", X"067A", X"0492", X"05AA", X"04EB", X"02A5", X"01BF", X"FEDC", X"FB44", X"F642", X"F4C3", X"F722", X"FDAA", X"001C", X"0210", X"024A", X"03B5", X"000F", X"FF5E", X"FE72", X"FE8F", X"FD6F", X"FC12", X"FA45", X"F977", X"FAAE", X"FE1F", X"043A", X"06E1", X"0578", X"0382", X"03E7", X"022C", X"01B6", X"013D", X"FE17", X"F71A", X"F2D8", X"F952", X"F9A0", X"FFFB", X"01A1", X"0037", X"015B", X"05B6", X"0270", X"FE8F", X"FC78", X"FBFC", X"FCD3", X"FD06", X"FEA4", X"0074", X"FD2D", X"FD72", X"029F", X"057B", X"04CC", X"0497", X"00CE", X"02E6", X"0180", X"FFBA", X"FCDC", X"F86F", X"F071", X"F820", X"FA45", X"01D1", X"009F", X"02B4", X"02E5", X"01E8", X"0280", X"FD25", X"FE56", X"FE32", X"00DE", X"02A4", X"02A0", X"FFDB", X"FFA5", X"FFBE", X"052F", X"05EC", X"0261", X"046B", X"028E", X"0249", X"0090", X"FDF5", X"FCD1", X"F81E", X"F33A", X"F952", X"FBBF", X"0260", X"015F", X"00C1", X"0159", X"01EC", X"0451", X"0142", X"0293", X"03DD", X"04D9", X"029E", X"03AF", X"FFDB", X"FC69", X"0079", X"0415", X"03C9", X"04D9", X"0654", X"051E", X"0130", X"00AD", X"FED2", X"FC59", X"F76C", X"F3DA", X"F9B7", X"FBEC", X"FBE3", X"FDC4", X"02AF", X"016C", X"02B8", X"07EB", X"04E2", X"073E", X"06C6", X"0589", X"02BB", X"FE9F", X"FD0D", X"FED7", X"00BC", X"02C6", X"03AD", X"035F", X"0497", X"0424", X"026E", X"035E", X"018D", X"FF8D", X"FB95", X"F809", X"F9F1", X"FD32", X"FEA7", X"FE57", X"02A7", X"0352", X"026F", X"06E1", X"0909", X"08A9", X"05A7", X"01B7", X"FEF9", X"FE36", X"FDC7", X"FE69", X"FEC0", X"02A8", X"02CE", X"041C", X"0547", X"030D", X"0359", X"0431", X"016A", X"019D", X"FD98", X"F5BC", X"F966", X"FEB2", X"FFDD", X"FF60", X"02E3", X"0413", X"FFFB", X"084E", X"0809", X"05DF", X"0452", X"00AF", X"FBA1", X"FC59", X"FD22", X"FBAF", X"FDB8", X"027A", X"0119", X"0230", X"035E", X"042D", X"02A0", X"032F", X"0331", X"018C", X"FD49", X"F81D", X"F583", X"FBCC", X"FE36", X"FFB8", X"017B", X"02FF", X"0344", X"0719", X"047C", X"030E", X"00A7", X"FFAB", X"FCEE", X"FC11", X"FBEE", X"FADB", X"FE60", X"0102", X"0204", X"0104", X"021B", X"0364", X"0095", X"FEB2", X"014F", X"0057", X"FCB8", X"F60B", X"F674", X"FDE0", X"FCDC", X"0374", X"00EE", X"02CD", X"0382", X"04E2", X"05CB", X"00D9", X"FEBB", X"FE24", X"FDF3", X"FC36", X"FB23", X"F852", X"FC1D", X"000D", X"00E5", X"FFC5", X"FFAA", X"FF89", X"003C", X"0083", X"01C8", X"FF05", X"FADB", X"F350", X"F861", X"0127", X"0201", X"FF9A", X"0220", X"FFDB", X"03F5", X"04E9", X"04A4", X"0097", X"FF65", X"FDBC", X"FB85", X"FB10", X"FAF7", X"F8D8", X"FE12", X"FEBC", X"0059", X"FF84", X"FF22", X"FF1C", X"0018", X"0032", X"FFD8", X"FD1E", X"F88E", X"F3A2", X"FB0B", X"FF7D", X"026C", X"FFA6", X"006C", X"FE73", X"00E5", X"0445", X"0000", X"00F9", X"00A3", X"FE12", X"FC87", X"FA69", X"FB0C", X"F968", X"FC8A", X"00C6", X"0025", X"FFEC", X"00AC", X"FF5D", X"FF75", X"FFD5", X"FDBB", X"FAD3", X"F7A7", X"F836", X"FF98", X"0035", X"0143", X"0051", X"FE90", X"FF93", X"FEE5", X"0435", X"0274", X"0095", X"FFF3", X"FF30", X"FC62", X"FC21", X"FA9C", X"FC5D", X"FC34", X"FE18", X"FF79", X"01E6", X"FF62", X"FF16", X"009C", X"FDD3", X"FE54", X"F95C", X"F933", X"FAA4", X"FF65", X"FC92", X"FF61", X"FF59", X"0034", X"0197", X"FE1C", X"018C", X"01B6", X"0279", X"02F0", X"FE1E", X"FED8", X"FDF9", X"FE57", X"FB97", X"FAF7", X"FD9B", X"006F", X"FF18", X"004B", X"FEC6", X"FFEA", X"FEAF", X"FD47", X"FBD4", X"FB17", X"FAE7", X"FF2F", X"0178", X"0144", X"0098", X"0111", X"FEA9", X"005C", X"02BC", X"0432", X"04F9", X"0272", X"0072", X"FF16", X"FE31", X"FE4D", X"FC16", X"FDE6", X"FD11", X"FEC4", X"FD6B", X"0127", X"0236", X"0206", X"FE7F", X"FDAB", X"FC92", X"FCA9", X"FE77", X"FFE9", X"0277", X"00AC", X"01FE", X"FF9F", X"00F1", X"053E", X"0813", X"080D", X"08FF", X"07D0", X"042E", X"032D", X"01A4", X"FF9F", X"FDDB", X"FE6B", X"FEF3", X"FE21", X"0192", X"014E", X"0191", X"024D", X"0367", X"0397", X"FE86", X"FFF5", X"FA2E", X"FCBC", X"FE33", X"FF9D", X"FE94", X"0020", X"FFB2", X"FFB9", X"04DB", X"0873", X"05DE", X"0670", X"09BF", X"0808", X"040B", X"0341", X"01C2", X"FF2B", X"0106", X"FF17", X"000E", X"0224", X"032C", X"0583", X"0603", X"0376", X"01FA", X"FD98", X"FEC4", X"FF23", X"FE16", X"006D", X"011C", X"0098", X"0158", X"005F", X"00F4", X"038A", X"079D", X"06D9", X"06E9", X"0621", X"032D", X"018E", X"FEFF", X"021D", X"054B", X"03DC", X"0652", X"045E", X"05AA", X"0503", X"0473", X"02B1", X"009B", X"FFA1", X"FFEC", X"FFDB", X"FED1", X"FF57", X"0177", X"FF84", X"FF24", X"013D", X"FEDE", X"0035", X"01D5", X"0103", X"01FE", X"0018", X"0242", X"FF19", X"016D", X"032F", X"0323", X"021E", X"0258", X"0105", X"031A", X"0195", X"0399", X"0289", X"0171", X"014E", X"0020", X"0055", X"FF89", X"0110"),
        (X"FEB6", X"00C4", X"0121", X"00D1", X"0111", X"004B", X"00B1", X"FF2D", X"00E2", X"FFC7", X"FFEA", X"FEEA", X"021A", X"FFDB", X"FFCF", X"01AD", X"0103", X"FE88", X"017B", X"FF58", X"00F4", X"008F", X"00C5", X"010B", X"FF5D", X"0036", X"00B1", X"FE1F", X"008E", X"00F7", X"FFCE", X"00F7", X"0014", X"FFB6", X"000B", X"FE56", X"FF7F", X"0106", X"0134", X"00AC", X"0214", X"0070", X"034A", X"0179", X"FFAF", X"01D0", X"0377", X"0193", X"028E", X"FF26", X"0034", X"FDA2", X"004A", X"0088", X"003A", X"028A", X"FFDC", X"0020", X"FF38", X"FDDE", X"FF71", X"00F8", X"000F", X"0003", X"00A4", X"01C7", X"0190", X"01F2", X"034C", X"0237", X"043A", X"0362", X"02F6", X"01EB", X"0137", X"0366", X"01EF", X"01B1", X"0307", X"FE24", X"FFDD", X"FE8D", X"FF87", X"00AE", X"001D", X"00C8", X"004A", X"FEFB", X"FF60", X"0072", X"0066", X"0166", X"03B1", X"06DF", X"05D2", X"0650", X"050B", X"03A8", X"0677", X"0679", X"0523", X"05C5", X"0238", X"0649", X"0639", X"0657", X"03E8", X"0257", X"019D", X"FE2D", X"004D", X"FEA6", X"FECE", X"0077", X"FF62", X"FDD5", X"00EA", X"0548", X"0595", X"07CD", X"08A6", X"0A17", X"0942", X"0BAD", X"0CC7", X"0DEF", X"0FC0", X"1166", X"0FDB", X"1077", X"0DC6", X"0C1B", X"0F8F", X"08C8", X"0AA1", X"05CB", X"0249", X"0097", X"022B", X"FF49", X"002A", X"0170", X"FF5F", X"01E9", X"04EF", X"0632", X"0801", X"0686", X"070A", X"076B", X"0743", X"066B", X"071E", X"0877", X"0C09", X"0CB4", X"0D83", X"090C", X"0616", X"028D", X"056A", X"065E", X"08E3", X"0C64", X"08B4", X"061D", X"0305", X"0121", X"FF16", X"FF91", X"FE70", X"FE6B", X"0290", X"066E", X"02E5", X"0468", X"03C8", X"0493", X"0401", X"FE97", X"00EC", X"004C", X"FF51", X"FE6E", X"FDF2", X"FF04", X"FD78", X"FF55", X"FF53", X"FF26", X"0465", X"09A5", X"0A18", X"057D", X"0525", X"01B4", X"013B", X"FFD9", X"FC80", X"FD94", X"0678", X"0670", X"010E", X"0217", X"021E", X"FEF6", X"FDA6", X"FECD", X"FB64", X"F982", X"F97B", X"F84B", X"F8A4", X"FA13", X"FC43", X"FF31", X"FFD0", X"00C6", X"042B", X"07AE", X"095A", X"0786", X"07A4", X"0168", X"00C8", X"FC39", X"0026", X"0215", X"041D", X"02D8", X"FEC4", X"FF1E", X"002B", X"FFB7", X"0076", X"FDCC", X"FD1C", X"FB21", X"FAA8", X"FA00", X"FDBF", X"FD23", X"FFF9", X"01B5", X"0010", X"01C7", X"00FB", X"03FD", X"047E", X"0A15", X"06E8", X"025A", X"FF71", X"FBDD", X"0185", X"FFC9", X"0298", X"014B", X"FC9D", X"FDBE", X"FE95", X"FDF0", X"FDCD", X"FD85", X"FB56", X"FB2E", X"F7C6", X"F94D", X"FEFA", X"0055", X"00D0", X"01C6", X"00AF", X"0225", X"0153", X"02A0", X"027D", X"05AA", X"035A", X"FDAD", X"0068", X"FD74", X"FE12", X"FEE0", X"04D4", X"FE9F", X"FB3F", X"FDE4", X"FF54", X"FCC4", X"FC17", X"FA76", X"FA37", X"F941", X"F8A8", X"FC24", X"FCA1", X"FEFC", X"FE11", X"FF44", X"FD9C", X"FD13", X"FEF5", X"FF4A", X"0264", X"0175", X"01D0", X"FF80", X"00BA", X"FDEE", X"FB84", X"FCD7", X"FDEC", X"FCD3", X"FCF3", X"FC9F", X"FEAD", X"FCD7", X"FD99", X"FCAB", X"FF60", X"FC0D", X"FAA1", X"F964", X"FC15", X"FD65", X"FC93", X"FCD9", X"FBA8", X"FAFA", X"FC32", X"FF0A", X"0095", X"00F0", X"02A3", X"00DA", X"FE9E", X"FE25", X"FD34", X"FC80", X"FBDB", X"FCFF", X"FF2E", X"FDC3", X"FE60", X"FF37", X"0161", X"018C", X"0497", X"0398", X"FC9F", X"FC53", X"FB74", X"FA3F", X"FC0F", X"FE45", X"FC62", X"FE87", X"FEBD", X"FE4E", X"04A7", X"FD16", X"FF58", X"FCFC", X"00A4", X"FF0F", X"FC94", X"FAFC", X"FAA7", X"FD8E", X"FE30", X"0064", X"0164", X"0341", X"02AB", X"08AC", X"0877", X"0346", X"FFF0", X"FE8E", X"FD03", X"FDCA", X"FE11", X"FE3A", X"0025", X"FE1E", X"0190", X"01EA", X"00B9", X"FD71", X"FCCB", X"FBD7", X"013F", X"FEA2", X"FD18", X"FCFE", X"FD06", X"FD59", X"001D", X"017C", X"0224", X"0387", X"0412", X"0545", X"05F4", X"0409", X"03A1", X"00AE", X"FF92", X"FF48", X"FEEE", X"FFA2", X"FEC3", X"FF44", X"0053", X"FF10", X"FFD8", X"FBA0", X"F6B9", X"FDF4", X"0245", X"FFC3", X"03AC", X"015B", X"FD45", X"FFBB", X"FE93", X"026B", X"0446", X"039B", X"0153", X"024A", X"0490", X"03C6", X"0688", X"02E2", X"FEB7", X"FD9B", X"FD82", X"FF48", X"FE28", X"FDFE", X"FD51", X"FF68", X"FC39", X"FA9C", X"FB4E", X"FD5F", X"FECB", X"0000", X"03F5", X"FF62", X"FABA", X"FCF1", X"FEAE", X"FE72", X"012F", X"0164", X"FFEA", X"006A", X"01B1", X"04E2", X"047A", X"01B7", X"FF35", X"FE2D", X"FD33", X"FD2D", X"FC85", X"0029", X"FE75", X"0000", X"FE84", X"FCD4", X"F9BD", X"FA98", X"00C8", X"FE91", X"0146", X"FEA7", X"FCAD", X"FF0E", X"FF1F", X"FF7C", X"FBEE", X"FDEC", X"FDB4", X"FF80", X"00E1", X"0162", X"0239", X"0071", X"FFFF", X"FE9F", X"FE05", X"FEF2", X"FEDF", X"010C", X"FFDE", X"FED1", X"FE73", X"F876", X"FCA9", X"FD4A", X"FE2B", X"0192", X"0093", X"FF23", X"FD6D", X"FF51", X"0038", X"FF71", X"FE7E", X"FCE3", X"FD5D", X"FEBE", X"01C4", X"001C", X"FF1F", X"0035", X"0190", X"FF35", X"FEE6", X"FE92", X"0085", X"0085", X"0024", X"0142", X"FD9F", X"F8E8", X"FC2B", X"FDBF", X"FFEA", X"FDBF", X"0049", X"019A", X"0037", X"0206", X"0500", X"0313", X"FFD8", X"FFE9", X"FF4B", X"006F", X"0108", X"01B6", X"00A3", X"02DF", X"0304", X"013B", X"0363", X"0145", X"0194", X"03D8", X"022D", X"00EE", X"FE65", X"F94E", X"FDF0", X"FED2", X"00CE", X"0213", X"04AB", X"0448", X"01D7", X"0472", X"098E", X"06ED", X"0446", X"044F", X"0443", X"04E0", X"02FB", X"00EE", X"0414", X"0501", X"02F8", X"0549", X"0530", X"02E4", X"0620", X"058F", X"05D1", X"0185", X"FB17", X"FB00", X"FE7C", X"000C", X"0039", X"0122", X"0567", X"0700", X"0190", X"067B", X"0913", X"08AE", X"06E5", X"05E1", X"0719", X"0663", X"0340", X"0340", X"0490", X"054D", X"02B9", X"07A6", X"071A", X"053F", X"050B", X"06D8", X"038C", X"0219", X"FDB7", X"FBE6", X"023C", X"00D3", X"FFF1", X"FFB9", X"056A", X"0581", X"0418", X"0489", X"07EE", X"0523", X"0483", X"065F", X"04E2", X"055D", X"03D2", X"0425", X"04B5", X"0531", X"0480", X"0789", X"07C6", X"07BE", X"0556", X"0639", X"02D9", X"FF53", X"FCAF", X"FEB6", X"0314", X"FFF7", X"0027", X"FE80", X"05A5", X"04AB", X"0091", X"FF56", X"0058", X"005D", X"0221", X"0484", X"0448", X"0549", X"050D", X"042C", X"0560", X"05E0", X"04C6", X"05E4", X"067C", X"069C", X"04F6", X"049C", X"017B", X"FF59", X"FCCF", X"FD8E", X"037A", X"FE9D", X"FF12", X"00D0", X"FE1D", X"0134", X"F8D9", X"F6A0", X"F78D", X"F919", X"FCC7", X"FFA8", X"0005", X"022A", X"02B5", X"032A", X"039F", X"014F", X"0390", X"011F", X"0229", X"0259", X"FF99", X"FCC6", X"FE92", X"FD1C", X"003B", X"0171", X"00B0", X"FD9F", X"0088", X"0136", X"FEDF", X"FF6C", X"F92B", X"F47D", X"F61D", X"F6BE", X"F739", X"F94E", X"FE6F", X"FCDA", X"FCC9", X"FEDF", X"FF6E", X"FF5D", X"FE69", X"FC72", X"FD90", X"FC30", X"FAC8", X"FAD6", X"FD39", X"FEC6", X"0192", X"FF3E", X"014A", X"0042", X"002A", X"0008", X"00C2", X"FF3A", X"FC34", X"F827", X"F5E4", X"F685", X"F673", X"F5FA", X"F60B", X"F87C", X"F91A", X"F745", X"F343", X"F5B5", X"FA54", X"F919", X"F7F6", X"F8DD", X"F8E4", X"FB5D", X"FD3E", X"FF27", X"0020", X"FFBE", X"0129", X"FF02", X"003A", X"010F", X"0073", X"FF0F", X"0098", X"FFCB", X"FD31", X"FD8B", X"FCE3", X"FC77", X"FBE2", X"FD11", X"FD31", X"FB53", X"F84F", X"FBEA", X"FBA1", X"FBAA", X"FAFC", X"FB86", X"FF94", X"FD28", X"FBCE", X"FE58", X"FFE9", X"FFE8", X"FE3A", X"0076")
);
    
    signal b1 : WORD_ARRAY(0 to unit_num1 - 1) := (	
	   (X"0124", X"FFFB", X"09CD", X"07F3", X"03BB", X"0388", X"FE1D", X"01DA", X"FDC4", X"059B", X"029C", X"FF6C", X"021D", X"F782", X"03A3", X"FC20", X"0071", X"FE04", X"FC08", X"FC62", X"FC13", X"FC73", X"FAFF", X"05F7", X"029C", X"FF68", X"08D3", X"0010", X"0477", X"013E", X"08E3", X"0B51", X"F66D", X"FC1C", X"F9F7", X"01AB", X"03E4", X"0597", X"FB0D", X"F955", X"0353", X"0538", X"0BE9", X"00C1", X"0203", X"FFDD", X"01D7", X"05FE", X"04AA", X"0193")
    );
    
    signal W2 : WORD_MAT(0 to unit_num2-1, 0 to input_dim2-1) := (	
        (X"F2FF", X"F7D0", X"F54B", X"F4A4", X"F1A6", X"F2EB", X"FFFC", X"F1D5", X"FB59", X"0604", X"022C", X"FFEB", X"F58D", X"F2D4", X"F5FF", X"00A3", X"F68D", X"F37E", X"F9B3", X"F207", X"FA44", X"FD23", X"086D", X"F274", X"0729", X"F86C", X"02F0", X"0887", X"F1A3", X"FBA0", X"039B", X"F50C", X"F65D", X"F2AF", X"02CA", X"0A3B", X"FF52", X"F71A", X"F2F9", X"F2BA", X"F612", X"0D79", X"EE6D", X"0036", X"F47A", X"F079", X"07E9", X"04BF", X"F829", X"FB1B"),
        (X"0345", X"F167", X"06EC", X"028F", X"06AC", X"0AF6", X"F321", X"05B8", X"F1F4", X"F75B", X"FA4E", X"F41F", X"F5F3", X"F5E0", X"06C0", X"F245", X"F7FC", X"FBEF", X"F0AE", X"05BB", X"02E0", X"F929", X"FE92", X"094B", X"F8B5", X"F0E7", X"F737", X"F701", X"FCCA", X"04D8", X"FEFA", X"F45E", X"018B", X"F1CB", X"F4AA", X"08B3", X"F969", X"FB1E", X"FA19", X"F39B", X"0264", X"0182", X"F800", X"F307", X"0909", X"018D", X"F3EA", X"F74D", X"FF93", X"FD08"),
        (X"F5EC", X"0BDB", X"F6D5", X"F450", X"F5C4", X"F596", X"FB0B", X"F124", X"0012", X"F908", X"0056", X"038F", X"05F9", X"F307", X"F931", X"F183", X"FDE7", X"EDB5", X"F4EB", X"08FD", X"FDA7", X"F174", X"0206", X"08A4", X"F83C", X"FBFC", X"F567", X"0B9F", X"FF26", X"F4D4", X"F35A", X"F932", X"F6A5", X"06EC", X"F9ED", X"069A", X"EEEC", X"F7FC", X"094F", X"068F", X"093B", X"F482", X"F596", X"044F", X"036C", X"038A", X"F818", X"F66C", X"F1B9", X"F884"),
        (X"F086", X"F29E", X"F6EA", X"F9D5", X"F4DC", X"04D7", X"FFBD", X"070B", X"0013", X"074F", X"EE76", X"0101", X"F5FB", X"094C", X"F3FD", X"015E", X"F1A3", X"044B", X"FEA9", X"F534", X"FBB4", X"FC04", X"F1A9", X"07C0", X"F243", X"FE3E", X"F53D", X"F21B", X"FBBC", X"F4AC", X"F808", X"F485", X"FC36", X"FA78", X"0375", X"F0FE", X"F032", X"F82E", X"03A7", X"F58A", X"0691", X"F52B", X"F5E8", X"047D", X"08C2", X"075A", X"F45B", X"04DE", X"07EF", X"F898"),
        (X"F797", X"FDDD", X"0BDF", X"FFEF", X"039A", X"F28B", X"00C8", X"F5E9", X"EFC9", X"F3D1", X"F28C", X"F928", X"0875", X"0576", X"03F1", X"036B", X"0052", X"FBDD", X"FA3E", X"F968", X"EF2A", X"F155", X"F60D", X"F735", X"0A9F", X"F7E6", X"024B", X"0492", X"F383", X"001F", X"F0B5", X"0973", X"F45D", X"FF54", X"F435", X"F6FF", X"F7DA", X"0910", X"F85F", X"02BA", X"F73E", X"F185", X"0409", X"F63B", X"F6F1", X"F239", X"EFDC", X"F4C4", X"FEEE", X"0351"),
        (X"094F", X"F3BC", X"0078", X"F537", X"00E4", X"FE83", X"EADD", X"0A2B", X"02C2", X"0E72", X"F3E8", X"0100", X"F97A", X"FCEE", X"EF07", X"F7E9", X"0106", X"FA9B", X"F1ED", X"FA35", X"F6AD", X"F765", X"EF9C", X"0620", X"0753", X"FCD4", X"074B", X"F41B", X"010C", X"01F1", X"07AC", X"0AB4", X"F0B6", X"F1FA", X"010C", X"F35A", X"FCBA", X"F55C", X"F468", X"F395", X"F59B", X"F3C5", X"0AF4", X"0459", X"F75B", X"F8BA", X"07D6", X"0290", X"F257", X"FB8C"),
        (X"0220", X"FAF5", X"0839", X"059F", X"F0D1", X"0BEB", X"EE63", X"FBA2", X"01C8", X"FB0C", X"015F", X"F2D4", X"0579", X"F7AF", X"F2C8", X"F233", X"FE29", X"F8E4", X"002E", X"F85C", X"F353", X"F325", X"082C", X"F015", X"F49A", X"FB81", X"062D", X"04F3", X"F17F", X"F86D", X"0305", X"F1DD", X"F5DE", X"FC5F", X"F477", X"089D", X"00A8", X"F350", X"F5C6", X"0049", X"EE99", X"FE9B", X"03EA", X"F171", X"F27D", X"08D8", X"F350", X"F341", X"F0E1", X"FF28"),
        (X"F273", X"07A8", X"F8CF", X"024D", X"0364", X"F712", X"FFAF", X"F034", X"F6C0", X"F8D7", X"05AF", X"F41D", X"F1A3", X"F323", X"0724", X"FE46", X"F37C", X"F676", X"FAD6", X"02AA", X"F358", X"FCBF", X"F4DF", X"F93A", X"F879", X"FB38", X"097D", X"F0E7", X"F8B6", X"F524", X"FB63", X"0821", X"0427", X"0043", X"EFEA", X"F293", X"F02E", X"0CC7", X"FA2B", X"F232", X"043F", X"0A4E", X"FBAF", X"FBED", X"09D4", X"FA22", X"FF37", X"0BF8", X"03D7", X"F216"),
        (X"056C", X"F9D7", X"F5DF", X"EEAE", X"010B", X"F4D6", X"F938", X"02B2", X"0227", X"EE4D", X"0186", X"FA83", X"EE70", X"0475", X"F68B", X"003E", X"0026", X"07DF", X"0075", X"08A9", X"FED7", X"0310", X"01C9", X"ED93", X"FD1B", X"FD81", X"F2B2", X"F1D5", X"FAB4", X"03C5", X"EE34", X"EE1F", X"0528", X"FB43", X"FB55", X"F2C9", X"0240", X"EAB1", X"09E0", X"FFE8", X"F20F", X"F2D7", X"F238", X"FAF5", X"F47E", X"F6DC", X"FB29", X"F4CB", X"F13D", X"FDFE"),
        (X"FF74", X"F79B", X"ECE5", X"FEE4", X"FBD9", X"F426", X"FE4A", X"F7D9", X"F2E3", X"F86B", X"F15E", X"FADA", X"0596", X"0703", X"05A4", X"002C", X"FA43", X"FCC8", X"FAB1", X"EB8B", X"07D5", X"068F", X"F8A2", X"F322", X"F222", X"F931", X"EDE8", X"FB8A", X"01B7", X"F41F", X"FFFC", X"0678", X"0672", X"F854", X"05E6", X"F99A", X"0120", X"067F", X"F07B", X"00B0", X"F639", X"FD43", X"FF1D", X"F2BF", X"F2A8", X"F4E7", X"07C4", X"F368", X"0413", X"F12B")
    );
    
    signal b2 : WORD_ARRAY(0 to unit_num2-1) := (    
        (X"F7FC", X"F8CF", X"F983", X"F93C", X"F8BF", X"FAA8", X"F961", X"F91C", X"F804", X"F961")
    );
    
    signal a2 : WORD_ARRAY(0 to unit_num1-1);
    signal a3 : WORD_ARRAY(0 to unit_num2-1);


begin
    
   
   ffu1: entity work.feed_forward_unit(Structural)
               generic map(
                           unit_num => 50,
                           input_dim => 784
               )
               
               port map( 
                         input => X,
                         weights => W1,
                         bias => b1,
                         a => a2
               );
               
               
  ffu2: entity work.feed_forward_unit(Structural)
                       generic map(
                                   unit_num => 10,
                                   input_dim => 50
                       )
                       
                       port map( 
                                 input => a2,
                                 weights => W2,
                                 bias => b2,
                                 a => a3
                       );



end Stimulus;
